//megafunction wizard: %Altera SOPC Builder%
//GENERATION: STANDARD
//VERSION: WM1.0


//Legal Notice: (C)2014 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module clocks_0_avalon_clocks_slave_arbitrator (
                                                 // inputs:
                                                  clk,
                                                  clocks_0_avalon_clocks_slave_readdata,
                                                  nios_system_clock_10_out_address_to_slave,
                                                  nios_system_clock_10_out_read,
                                                  nios_system_clock_10_out_write,
                                                  nios_system_clock_11_out_address_to_slave,
                                                  nios_system_clock_11_out_read,
                                                  nios_system_clock_11_out_write,
                                                  nios_system_clock_8_out_address_to_slave,
                                                  nios_system_clock_8_out_read,
                                                  nios_system_clock_8_out_write,
                                                  nios_system_clock_9_out_address_to_slave,
                                                  nios_system_clock_9_out_read,
                                                  nios_system_clock_9_out_write,
                                                  reset_n,

                                                 // outputs:
                                                  clocks_0_avalon_clocks_slave_address,
                                                  clocks_0_avalon_clocks_slave_readdata_from_sa,
                                                  d1_clocks_0_avalon_clocks_slave_end_xfer,
                                                  nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave,
                                                  nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave
                                               )
;

  output           clocks_0_avalon_clocks_slave_address;
  output  [  7: 0] clocks_0_avalon_clocks_slave_readdata_from_sa;
  output           d1_clocks_0_avalon_clocks_slave_end_xfer;
  output           nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave;
  output           nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave;
  input            clk;
  input   [  7: 0] clocks_0_avalon_clocks_slave_readdata;
  input            nios_system_clock_10_out_address_to_slave;
  input            nios_system_clock_10_out_read;
  input            nios_system_clock_10_out_write;
  input            nios_system_clock_11_out_address_to_slave;
  input            nios_system_clock_11_out_read;
  input            nios_system_clock_11_out_write;
  input            nios_system_clock_8_out_address_to_slave;
  input            nios_system_clock_8_out_read;
  input            nios_system_clock_8_out_write;
  input            nios_system_clock_9_out_address_to_slave;
  input            nios_system_clock_9_out_read;
  input            nios_system_clock_9_out_write;
  input            reset_n;

  wire             clocks_0_avalon_clocks_slave_address;
  wire             clocks_0_avalon_clocks_slave_allgrants;
  wire             clocks_0_avalon_clocks_slave_allow_new_arb_cycle;
  wire             clocks_0_avalon_clocks_slave_any_bursting_master_saved_grant;
  wire             clocks_0_avalon_clocks_slave_any_continuerequest;
  reg     [  3: 0] clocks_0_avalon_clocks_slave_arb_addend;
  wire             clocks_0_avalon_clocks_slave_arb_counter_enable;
  reg              clocks_0_avalon_clocks_slave_arb_share_counter;
  wire             clocks_0_avalon_clocks_slave_arb_share_counter_next_value;
  wire             clocks_0_avalon_clocks_slave_arb_share_set_values;
  wire    [  3: 0] clocks_0_avalon_clocks_slave_arb_winner;
  wire             clocks_0_avalon_clocks_slave_arbitration_holdoff_internal;
  wire             clocks_0_avalon_clocks_slave_beginbursttransfer_internal;
  wire             clocks_0_avalon_clocks_slave_begins_xfer;
  wire    [  7: 0] clocks_0_avalon_clocks_slave_chosen_master_double_vector;
  wire    [  3: 0] clocks_0_avalon_clocks_slave_chosen_master_rot_left;
  wire             clocks_0_avalon_clocks_slave_end_xfer;
  wire             clocks_0_avalon_clocks_slave_firsttransfer;
  wire    [  3: 0] clocks_0_avalon_clocks_slave_grant_vector;
  wire             clocks_0_avalon_clocks_slave_in_a_read_cycle;
  wire             clocks_0_avalon_clocks_slave_in_a_write_cycle;
  wire    [  3: 0] clocks_0_avalon_clocks_slave_master_qreq_vector;
  wire             clocks_0_avalon_clocks_slave_non_bursting_master_requests;
  wire    [  7: 0] clocks_0_avalon_clocks_slave_readdata_from_sa;
  reg              clocks_0_avalon_clocks_slave_reg_firsttransfer;
  reg     [  3: 0] clocks_0_avalon_clocks_slave_saved_chosen_master_vector;
  reg              clocks_0_avalon_clocks_slave_slavearbiterlockenable;
  wire             clocks_0_avalon_clocks_slave_slavearbiterlockenable2;
  wire             clocks_0_avalon_clocks_slave_unreg_firsttransfer;
  wire             clocks_0_avalon_clocks_slave_waits_for_read;
  wire             clocks_0_avalon_clocks_slave_waits_for_write;
  reg              d1_clocks_0_avalon_clocks_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_clocks_0_avalon_clocks_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_nios_system_clock_10_out_granted_slave_clocks_0_avalon_clocks_slave;
  reg              last_cycle_nios_system_clock_11_out_granted_slave_clocks_0_avalon_clocks_slave;
  reg              last_cycle_nios_system_clock_8_out_granted_slave_clocks_0_avalon_clocks_slave;
  reg              last_cycle_nios_system_clock_9_out_granted_slave_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_10_out_arbiterlock;
  wire             nios_system_clock_10_out_arbiterlock2;
  wire             nios_system_clock_10_out_continuerequest;
  wire             nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave;
  reg              nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
  wire             nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in;
  wire             nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_10_out_saved_grant_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_11_out_arbiterlock;
  wire             nios_system_clock_11_out_arbiterlock2;
  wire             nios_system_clock_11_out_continuerequest;
  wire             nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave;
  reg              nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
  wire             nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in;
  wire             nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_11_out_saved_grant_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_8_out_arbiterlock;
  wire             nios_system_clock_8_out_arbiterlock2;
  wire             nios_system_clock_8_out_continuerequest;
  wire             nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave;
  reg              nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
  wire             nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in;
  wire             nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_8_out_saved_grant_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_9_out_arbiterlock;
  wire             nios_system_clock_9_out_arbiterlock2;
  wire             nios_system_clock_9_out_continuerequest;
  wire             nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave;
  reg              nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
  wire             nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in;
  wire             nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_9_out_saved_grant_clocks_0_avalon_clocks_slave;
  wire             p1_nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
  wire             p1_nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
  wire             p1_nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
  wire             p1_nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
  wire             wait_for_clocks_0_avalon_clocks_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~clocks_0_avalon_clocks_slave_end_xfer;
    end


  assign clocks_0_avalon_clocks_slave_begins_xfer = ~d1_reasons_to_wait & ((nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave | nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave | nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave | nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave));
  //assign clocks_0_avalon_clocks_slave_readdata_from_sa = clocks_0_avalon_clocks_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign clocks_0_avalon_clocks_slave_readdata_from_sa = clocks_0_avalon_clocks_slave_readdata;

  assign nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave = ((1) & (nios_system_clock_10_out_read | nios_system_clock_10_out_write)) & nios_system_clock_10_out_read;
  //clocks_0_avalon_clocks_slave_arb_share_counter set values, which is an e_mux
  assign clocks_0_avalon_clocks_slave_arb_share_set_values = 1;

  //clocks_0_avalon_clocks_slave_non_bursting_master_requests mux, which is an e_mux
  assign clocks_0_avalon_clocks_slave_non_bursting_master_requests = nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave |
    nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave;

  //clocks_0_avalon_clocks_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign clocks_0_avalon_clocks_slave_any_bursting_master_saved_grant = 0;

  //clocks_0_avalon_clocks_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign clocks_0_avalon_clocks_slave_arb_share_counter_next_value = clocks_0_avalon_clocks_slave_firsttransfer ? (clocks_0_avalon_clocks_slave_arb_share_set_values - 1) : |clocks_0_avalon_clocks_slave_arb_share_counter ? (clocks_0_avalon_clocks_slave_arb_share_counter - 1) : 0;

  //clocks_0_avalon_clocks_slave_allgrants all slave grants, which is an e_mux
  assign clocks_0_avalon_clocks_slave_allgrants = (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector) |
    (|clocks_0_avalon_clocks_slave_grant_vector);

  //clocks_0_avalon_clocks_slave_end_xfer assignment, which is an e_assign
  assign clocks_0_avalon_clocks_slave_end_xfer = ~(clocks_0_avalon_clocks_slave_waits_for_read | clocks_0_avalon_clocks_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_clocks_0_avalon_clocks_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_clocks_0_avalon_clocks_slave = clocks_0_avalon_clocks_slave_end_xfer & (~clocks_0_avalon_clocks_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //clocks_0_avalon_clocks_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign clocks_0_avalon_clocks_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_clocks_0_avalon_clocks_slave & clocks_0_avalon_clocks_slave_allgrants) | (end_xfer_arb_share_counter_term_clocks_0_avalon_clocks_slave & ~clocks_0_avalon_clocks_slave_non_bursting_master_requests);

  //clocks_0_avalon_clocks_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clocks_0_avalon_clocks_slave_arb_share_counter <= 0;
      else if (clocks_0_avalon_clocks_slave_arb_counter_enable)
          clocks_0_avalon_clocks_slave_arb_share_counter <= clocks_0_avalon_clocks_slave_arb_share_counter_next_value;
    end


  //clocks_0_avalon_clocks_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clocks_0_avalon_clocks_slave_slavearbiterlockenable <= 0;
      else if ((|clocks_0_avalon_clocks_slave_master_qreq_vector & end_xfer_arb_share_counter_term_clocks_0_avalon_clocks_slave) | (end_xfer_arb_share_counter_term_clocks_0_avalon_clocks_slave & ~clocks_0_avalon_clocks_slave_non_bursting_master_requests))
          clocks_0_avalon_clocks_slave_slavearbiterlockenable <= |clocks_0_avalon_clocks_slave_arb_share_counter_next_value;
    end


  //nios_system_clock_10/out clocks_0/avalon_clocks_slave arbiterlock, which is an e_assign
  assign nios_system_clock_10_out_arbiterlock = clocks_0_avalon_clocks_slave_slavearbiterlockenable & nios_system_clock_10_out_continuerequest;

  //clocks_0_avalon_clocks_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign clocks_0_avalon_clocks_slave_slavearbiterlockenable2 = |clocks_0_avalon_clocks_slave_arb_share_counter_next_value;

  //nios_system_clock_10/out clocks_0/avalon_clocks_slave arbiterlock2, which is an e_assign
  assign nios_system_clock_10_out_arbiterlock2 = clocks_0_avalon_clocks_slave_slavearbiterlockenable2 & nios_system_clock_10_out_continuerequest;

  //nios_system_clock_11/out clocks_0/avalon_clocks_slave arbiterlock, which is an e_assign
  assign nios_system_clock_11_out_arbiterlock = clocks_0_avalon_clocks_slave_slavearbiterlockenable & nios_system_clock_11_out_continuerequest;

  //nios_system_clock_11/out clocks_0/avalon_clocks_slave arbiterlock2, which is an e_assign
  assign nios_system_clock_11_out_arbiterlock2 = clocks_0_avalon_clocks_slave_slavearbiterlockenable2 & nios_system_clock_11_out_continuerequest;

  //nios_system_clock_11/out granted clocks_0/avalon_clocks_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_11_out_granted_slave_clocks_0_avalon_clocks_slave <= 0;
      else 
        last_cycle_nios_system_clock_11_out_granted_slave_clocks_0_avalon_clocks_slave <= nios_system_clock_11_out_saved_grant_clocks_0_avalon_clocks_slave ? 1 : (clocks_0_avalon_clocks_slave_arbitration_holdoff_internal | ~nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave) ? 0 : last_cycle_nios_system_clock_11_out_granted_slave_clocks_0_avalon_clocks_slave;
    end


  //nios_system_clock_11_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_11_out_continuerequest = (last_cycle_nios_system_clock_11_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave) |
    (last_cycle_nios_system_clock_11_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave) |
    (last_cycle_nios_system_clock_11_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave);

  //clocks_0_avalon_clocks_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  assign clocks_0_avalon_clocks_slave_any_continuerequest = nios_system_clock_11_out_continuerequest |
    nios_system_clock_8_out_continuerequest |
    nios_system_clock_9_out_continuerequest |
    nios_system_clock_10_out_continuerequest |
    nios_system_clock_8_out_continuerequest |
    nios_system_clock_9_out_continuerequest |
    nios_system_clock_10_out_continuerequest |
    nios_system_clock_11_out_continuerequest |
    nios_system_clock_9_out_continuerequest |
    nios_system_clock_10_out_continuerequest |
    nios_system_clock_11_out_continuerequest |
    nios_system_clock_8_out_continuerequest;

  //nios_system_clock_8/out clocks_0/avalon_clocks_slave arbiterlock, which is an e_assign
  assign nios_system_clock_8_out_arbiterlock = clocks_0_avalon_clocks_slave_slavearbiterlockenable & nios_system_clock_8_out_continuerequest;

  //nios_system_clock_8/out clocks_0/avalon_clocks_slave arbiterlock2, which is an e_assign
  assign nios_system_clock_8_out_arbiterlock2 = clocks_0_avalon_clocks_slave_slavearbiterlockenable2 & nios_system_clock_8_out_continuerequest;

  //nios_system_clock_8/out granted clocks_0/avalon_clocks_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_8_out_granted_slave_clocks_0_avalon_clocks_slave <= 0;
      else 
        last_cycle_nios_system_clock_8_out_granted_slave_clocks_0_avalon_clocks_slave <= nios_system_clock_8_out_saved_grant_clocks_0_avalon_clocks_slave ? 1 : (clocks_0_avalon_clocks_slave_arbitration_holdoff_internal | ~nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave) ? 0 : last_cycle_nios_system_clock_8_out_granted_slave_clocks_0_avalon_clocks_slave;
    end


  //nios_system_clock_8_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_8_out_continuerequest = (last_cycle_nios_system_clock_8_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave) |
    (last_cycle_nios_system_clock_8_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave) |
    (last_cycle_nios_system_clock_8_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave);

  //nios_system_clock_9/out clocks_0/avalon_clocks_slave arbiterlock, which is an e_assign
  assign nios_system_clock_9_out_arbiterlock = clocks_0_avalon_clocks_slave_slavearbiterlockenable & nios_system_clock_9_out_continuerequest;

  //nios_system_clock_9/out clocks_0/avalon_clocks_slave arbiterlock2, which is an e_assign
  assign nios_system_clock_9_out_arbiterlock2 = clocks_0_avalon_clocks_slave_slavearbiterlockenable2 & nios_system_clock_9_out_continuerequest;

  //nios_system_clock_9/out granted clocks_0/avalon_clocks_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_9_out_granted_slave_clocks_0_avalon_clocks_slave <= 0;
      else 
        last_cycle_nios_system_clock_9_out_granted_slave_clocks_0_avalon_clocks_slave <= nios_system_clock_9_out_saved_grant_clocks_0_avalon_clocks_slave ? 1 : (clocks_0_avalon_clocks_slave_arbitration_holdoff_internal | ~nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave) ? 0 : last_cycle_nios_system_clock_9_out_granted_slave_clocks_0_avalon_clocks_slave;
    end


  //nios_system_clock_9_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_9_out_continuerequest = (last_cycle_nios_system_clock_9_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave) |
    (last_cycle_nios_system_clock_9_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave) |
    (last_cycle_nios_system_clock_9_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave);

  assign nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave = nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave & ~((nios_system_clock_10_out_read & ((|nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register))) | nios_system_clock_11_out_arbiterlock | nios_system_clock_8_out_arbiterlock | nios_system_clock_9_out_arbiterlock);
  //nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in = nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_10_out_read & ~clocks_0_avalon_clocks_slave_waits_for_read & ~(|nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register);

  //shift register p1 nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register = {nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register, nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in};

  //nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register <= 0;
      else 
        nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register <= p1_nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
    end


  //local readdatavalid nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave, which is an e_mux
  assign nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave = nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;

  assign nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave = ((1) & (nios_system_clock_11_out_read | nios_system_clock_11_out_write)) & nios_system_clock_11_out_read;
  //nios_system_clock_10/out granted clocks_0/avalon_clocks_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_10_out_granted_slave_clocks_0_avalon_clocks_slave <= 0;
      else 
        last_cycle_nios_system_clock_10_out_granted_slave_clocks_0_avalon_clocks_slave <= nios_system_clock_10_out_saved_grant_clocks_0_avalon_clocks_slave ? 1 : (clocks_0_avalon_clocks_slave_arbitration_holdoff_internal | ~nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave) ? 0 : last_cycle_nios_system_clock_10_out_granted_slave_clocks_0_avalon_clocks_slave;
    end


  //nios_system_clock_10_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_10_out_continuerequest = (last_cycle_nios_system_clock_10_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave) |
    (last_cycle_nios_system_clock_10_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave) |
    (last_cycle_nios_system_clock_10_out_granted_slave_clocks_0_avalon_clocks_slave & nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave);

  assign nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave = nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave & ~((nios_system_clock_11_out_read & ((|nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register))) | nios_system_clock_10_out_arbiterlock | nios_system_clock_8_out_arbiterlock | nios_system_clock_9_out_arbiterlock);
  //nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in = nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_11_out_read & ~clocks_0_avalon_clocks_slave_waits_for_read & ~(|nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register);

  //shift register p1 nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register = {nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register, nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in};

  //nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register <= 0;
      else 
        nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register <= p1_nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
    end


  //local readdatavalid nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave, which is an e_mux
  assign nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave = nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;

  assign nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave = ((1) & (nios_system_clock_8_out_read | nios_system_clock_8_out_write)) & nios_system_clock_8_out_read;
  assign nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave = nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave & ~((nios_system_clock_8_out_read & ((|nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register))) | nios_system_clock_10_out_arbiterlock | nios_system_clock_11_out_arbiterlock | nios_system_clock_9_out_arbiterlock);
  //nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in = nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_8_out_read & ~clocks_0_avalon_clocks_slave_waits_for_read & ~(|nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register);

  //shift register p1 nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register = {nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register, nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in};

  //nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register <= 0;
      else 
        nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register <= p1_nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
    end


  //local readdatavalid nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave, which is an e_mux
  assign nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave = nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;

  assign nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave = ((1) & (nios_system_clock_9_out_read | nios_system_clock_9_out_write)) & nios_system_clock_9_out_read;
  assign nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave = nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave & ~((nios_system_clock_9_out_read & ((|nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register))) | nios_system_clock_10_out_arbiterlock | nios_system_clock_11_out_arbiterlock | nios_system_clock_8_out_arbiterlock);
  //nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in = nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_9_out_read & ~clocks_0_avalon_clocks_slave_waits_for_read & ~(|nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register);

  //shift register p1 nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register = {nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register, nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register_in};

  //nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register <= 0;
      else 
        nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register <= p1_nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;
    end


  //local readdatavalid nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave, which is an e_mux
  assign nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave = nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave_shift_register;

  //allow new arb cycle for clocks_0/avalon_clocks_slave, which is an e_assign
  assign clocks_0_avalon_clocks_slave_allow_new_arb_cycle = ~nios_system_clock_10_out_arbiterlock & ~nios_system_clock_11_out_arbiterlock & ~nios_system_clock_8_out_arbiterlock & ~nios_system_clock_9_out_arbiterlock;

  //nios_system_clock_9/out assignment into master qualified-requests vector for clocks_0/avalon_clocks_slave, which is an e_assign
  assign clocks_0_avalon_clocks_slave_master_qreq_vector[0] = nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave;

  //nios_system_clock_9/out grant clocks_0/avalon_clocks_slave, which is an e_assign
  assign nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave = clocks_0_avalon_clocks_slave_grant_vector[0];

  //nios_system_clock_9/out saved-grant clocks_0/avalon_clocks_slave, which is an e_assign
  assign nios_system_clock_9_out_saved_grant_clocks_0_avalon_clocks_slave = clocks_0_avalon_clocks_slave_arb_winner[0] && nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave;

  //nios_system_clock_8/out assignment into master qualified-requests vector for clocks_0/avalon_clocks_slave, which is an e_assign
  assign clocks_0_avalon_clocks_slave_master_qreq_vector[1] = nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave;

  //nios_system_clock_8/out grant clocks_0/avalon_clocks_slave, which is an e_assign
  assign nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave = clocks_0_avalon_clocks_slave_grant_vector[1];

  //nios_system_clock_8/out saved-grant clocks_0/avalon_clocks_slave, which is an e_assign
  assign nios_system_clock_8_out_saved_grant_clocks_0_avalon_clocks_slave = clocks_0_avalon_clocks_slave_arb_winner[1] && nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave;

  //nios_system_clock_11/out assignment into master qualified-requests vector for clocks_0/avalon_clocks_slave, which is an e_assign
  assign clocks_0_avalon_clocks_slave_master_qreq_vector[2] = nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave;

  //nios_system_clock_11/out grant clocks_0/avalon_clocks_slave, which is an e_assign
  assign nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave = clocks_0_avalon_clocks_slave_grant_vector[2];

  //nios_system_clock_11/out saved-grant clocks_0/avalon_clocks_slave, which is an e_assign
  assign nios_system_clock_11_out_saved_grant_clocks_0_avalon_clocks_slave = clocks_0_avalon_clocks_slave_arb_winner[2] && nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave;

  //nios_system_clock_10/out assignment into master qualified-requests vector for clocks_0/avalon_clocks_slave, which is an e_assign
  assign clocks_0_avalon_clocks_slave_master_qreq_vector[3] = nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave;

  //nios_system_clock_10/out grant clocks_0/avalon_clocks_slave, which is an e_assign
  assign nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave = clocks_0_avalon_clocks_slave_grant_vector[3];

  //nios_system_clock_10/out saved-grant clocks_0/avalon_clocks_slave, which is an e_assign
  assign nios_system_clock_10_out_saved_grant_clocks_0_avalon_clocks_slave = clocks_0_avalon_clocks_slave_arb_winner[3] && nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave;

  //clocks_0/avalon_clocks_slave chosen-master double-vector, which is an e_assign
  assign clocks_0_avalon_clocks_slave_chosen_master_double_vector = {clocks_0_avalon_clocks_slave_master_qreq_vector, clocks_0_avalon_clocks_slave_master_qreq_vector} & ({~clocks_0_avalon_clocks_slave_master_qreq_vector, ~clocks_0_avalon_clocks_slave_master_qreq_vector} + clocks_0_avalon_clocks_slave_arb_addend);

  //stable onehot encoding of arb winner
  assign clocks_0_avalon_clocks_slave_arb_winner = (clocks_0_avalon_clocks_slave_allow_new_arb_cycle & | clocks_0_avalon_clocks_slave_grant_vector) ? clocks_0_avalon_clocks_slave_grant_vector : clocks_0_avalon_clocks_slave_saved_chosen_master_vector;

  //saved clocks_0_avalon_clocks_slave_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clocks_0_avalon_clocks_slave_saved_chosen_master_vector <= 0;
      else if (clocks_0_avalon_clocks_slave_allow_new_arb_cycle)
          clocks_0_avalon_clocks_slave_saved_chosen_master_vector <= |clocks_0_avalon_clocks_slave_grant_vector ? clocks_0_avalon_clocks_slave_grant_vector : clocks_0_avalon_clocks_slave_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign clocks_0_avalon_clocks_slave_grant_vector = {(clocks_0_avalon_clocks_slave_chosen_master_double_vector[3] | clocks_0_avalon_clocks_slave_chosen_master_double_vector[7]),
    (clocks_0_avalon_clocks_slave_chosen_master_double_vector[2] | clocks_0_avalon_clocks_slave_chosen_master_double_vector[6]),
    (clocks_0_avalon_clocks_slave_chosen_master_double_vector[1] | clocks_0_avalon_clocks_slave_chosen_master_double_vector[5]),
    (clocks_0_avalon_clocks_slave_chosen_master_double_vector[0] | clocks_0_avalon_clocks_slave_chosen_master_double_vector[4])};

  //clocks_0/avalon_clocks_slave chosen master rotated left, which is an e_assign
  assign clocks_0_avalon_clocks_slave_chosen_master_rot_left = (clocks_0_avalon_clocks_slave_arb_winner << 1) ? (clocks_0_avalon_clocks_slave_arb_winner << 1) : 1;

  //clocks_0/avalon_clocks_slave's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clocks_0_avalon_clocks_slave_arb_addend <= 1;
      else if (|clocks_0_avalon_clocks_slave_grant_vector)
          clocks_0_avalon_clocks_slave_arb_addend <= clocks_0_avalon_clocks_slave_end_xfer? clocks_0_avalon_clocks_slave_chosen_master_rot_left : clocks_0_avalon_clocks_slave_grant_vector;
    end


  //clocks_0_avalon_clocks_slave_firsttransfer first transaction, which is an e_assign
  assign clocks_0_avalon_clocks_slave_firsttransfer = clocks_0_avalon_clocks_slave_begins_xfer ? clocks_0_avalon_clocks_slave_unreg_firsttransfer : clocks_0_avalon_clocks_slave_reg_firsttransfer;

  //clocks_0_avalon_clocks_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign clocks_0_avalon_clocks_slave_unreg_firsttransfer = ~(clocks_0_avalon_clocks_slave_slavearbiterlockenable & clocks_0_avalon_clocks_slave_any_continuerequest);

  //clocks_0_avalon_clocks_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          clocks_0_avalon_clocks_slave_reg_firsttransfer <= 1'b1;
      else if (clocks_0_avalon_clocks_slave_begins_xfer)
          clocks_0_avalon_clocks_slave_reg_firsttransfer <= clocks_0_avalon_clocks_slave_unreg_firsttransfer;
    end


  //clocks_0_avalon_clocks_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign clocks_0_avalon_clocks_slave_beginbursttransfer_internal = clocks_0_avalon_clocks_slave_begins_xfer;

  //clocks_0_avalon_clocks_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign clocks_0_avalon_clocks_slave_arbitration_holdoff_internal = clocks_0_avalon_clocks_slave_begins_xfer & clocks_0_avalon_clocks_slave_firsttransfer;

  //clocks_0_avalon_clocks_slave_address mux, which is an e_mux
  assign clocks_0_avalon_clocks_slave_address = (nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave)? nios_system_clock_10_out_address_to_slave :
    (nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave)? nios_system_clock_11_out_address_to_slave :
    (nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave)? nios_system_clock_8_out_address_to_slave :
    nios_system_clock_9_out_address_to_slave;

  //d1_clocks_0_avalon_clocks_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_clocks_0_avalon_clocks_slave_end_xfer <= 1;
      else 
        d1_clocks_0_avalon_clocks_slave_end_xfer <= clocks_0_avalon_clocks_slave_end_xfer;
    end


  //clocks_0_avalon_clocks_slave_waits_for_read in a cycle, which is an e_mux
  assign clocks_0_avalon_clocks_slave_waits_for_read = clocks_0_avalon_clocks_slave_in_a_read_cycle & 0;

  //clocks_0_avalon_clocks_slave_in_a_read_cycle assignment, which is an e_assign
  assign clocks_0_avalon_clocks_slave_in_a_read_cycle = (nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_10_out_read) | (nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_11_out_read) | (nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_8_out_read) | (nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_9_out_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = clocks_0_avalon_clocks_slave_in_a_read_cycle;

  //clocks_0_avalon_clocks_slave_waits_for_write in a cycle, which is an e_mux
  assign clocks_0_avalon_clocks_slave_waits_for_write = clocks_0_avalon_clocks_slave_in_a_write_cycle & 0;

  //clocks_0_avalon_clocks_slave_in_a_write_cycle assignment, which is an e_assign
  assign clocks_0_avalon_clocks_slave_in_a_write_cycle = (nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_10_out_write) | (nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_11_out_write) | (nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_8_out_write) | (nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave & nios_system_clock_9_out_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = clocks_0_avalon_clocks_slave_in_a_write_cycle;

  assign wait_for_clocks_0_avalon_clocks_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //clocks_0/avalon_clocks_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave + nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave + nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave + nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (nios_system_clock_10_out_saved_grant_clocks_0_avalon_clocks_slave + nios_system_clock_11_out_saved_grant_clocks_0_avalon_clocks_slave + nios_system_clock_8_out_saved_grant_clocks_0_avalon_clocks_slave + nios_system_clock_9_out_saved_grant_clocks_0_avalon_clocks_slave > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_0_jtag_debug_module_arbitrator (
                                            // inputs:
                                             clk,
                                             cpu_0_data_master_address_to_slave,
                                             cpu_0_data_master_byteenable,
                                             cpu_0_data_master_debugaccess,
                                             cpu_0_data_master_latency_counter,
                                             cpu_0_data_master_read,
                                             cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                             cpu_0_data_master_write,
                                             cpu_0_data_master_writedata,
                                             cpu_0_instruction_master_address_to_slave,
                                             cpu_0_instruction_master_latency_counter,
                                             cpu_0_instruction_master_read,
                                             cpu_0_jtag_debug_module_readdata,
                                             cpu_0_jtag_debug_module_resetrequest,
                                             reset_n,

                                            // outputs:
                                             cpu_0_data_master_granted_cpu_0_jtag_debug_module,
                                             cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module,
                                             cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module,
                                             cpu_0_data_master_requests_cpu_0_jtag_debug_module,
                                             cpu_0_instruction_master_granted_cpu_0_jtag_debug_module,
                                             cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module,
                                             cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module,
                                             cpu_0_instruction_master_requests_cpu_0_jtag_debug_module,
                                             cpu_0_jtag_debug_module_address,
                                             cpu_0_jtag_debug_module_begintransfer,
                                             cpu_0_jtag_debug_module_byteenable,
                                             cpu_0_jtag_debug_module_chipselect,
                                             cpu_0_jtag_debug_module_debugaccess,
                                             cpu_0_jtag_debug_module_readdata_from_sa,
                                             cpu_0_jtag_debug_module_resetrequest_from_sa,
                                             cpu_0_jtag_debug_module_write,
                                             cpu_0_jtag_debug_module_writedata,
                                             d1_cpu_0_jtag_debug_module_end_xfer
                                          )
;

  output           cpu_0_data_master_granted_cpu_0_jtag_debug_module;
  output           cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  output           cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module;
  output           cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  output           cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  output           cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  output           cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module;
  output           cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  output  [  8: 0] cpu_0_jtag_debug_module_address;
  output           cpu_0_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_0_jtag_debug_module_byteenable;
  output           cpu_0_jtag_debug_module_chipselect;
  output           cpu_0_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_0_jtag_debug_module_readdata_from_sa;
  output           cpu_0_jtag_debug_module_resetrequest_from_sa;
  output           cpu_0_jtag_debug_module_write;
  output  [ 31: 0] cpu_0_jtag_debug_module_writedata;
  output           d1_cpu_0_jtag_debug_module_end_xfer;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input            cpu_0_data_master_debugaccess;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input            cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input   [ 31: 0] cpu_0_jtag_debug_module_readdata;
  input            cpu_0_jtag_debug_module_resetrequest;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module;
  wire    [  8: 0] cpu_0_jtag_debug_module_address;
  wire             cpu_0_jtag_debug_module_allgrants;
  wire             cpu_0_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_0_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_0_jtag_debug_module_any_continuerequest;
  reg     [  1: 0] cpu_0_jtag_debug_module_arb_addend;
  wire             cpu_0_jtag_debug_module_arb_counter_enable;
  reg     [  2: 0] cpu_0_jtag_debug_module_arb_share_counter;
  wire    [  2: 0] cpu_0_jtag_debug_module_arb_share_counter_next_value;
  wire    [  2: 0] cpu_0_jtag_debug_module_arb_share_set_values;
  wire    [  1: 0] cpu_0_jtag_debug_module_arb_winner;
  wire             cpu_0_jtag_debug_module_arbitration_holdoff_internal;
  wire             cpu_0_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_0_jtag_debug_module_begins_xfer;
  wire             cpu_0_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_0_jtag_debug_module_byteenable;
  wire             cpu_0_jtag_debug_module_chipselect;
  wire    [  3: 0] cpu_0_jtag_debug_module_chosen_master_double_vector;
  wire    [  1: 0] cpu_0_jtag_debug_module_chosen_master_rot_left;
  wire             cpu_0_jtag_debug_module_debugaccess;
  wire             cpu_0_jtag_debug_module_end_xfer;
  wire             cpu_0_jtag_debug_module_firsttransfer;
  wire    [  1: 0] cpu_0_jtag_debug_module_grant_vector;
  wire             cpu_0_jtag_debug_module_in_a_read_cycle;
  wire             cpu_0_jtag_debug_module_in_a_write_cycle;
  wire    [  1: 0] cpu_0_jtag_debug_module_master_qreq_vector;
  wire             cpu_0_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_0_jtag_debug_module_readdata_from_sa;
  reg              cpu_0_jtag_debug_module_reg_firsttransfer;
  wire             cpu_0_jtag_debug_module_resetrequest_from_sa;
  reg     [  1: 0] cpu_0_jtag_debug_module_saved_chosen_master_vector;
  reg              cpu_0_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_0_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_0_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_0_jtag_debug_module_waits_for_read;
  wire             cpu_0_jtag_debug_module_waits_for_write;
  wire             cpu_0_jtag_debug_module_write;
  wire    [ 31: 0] cpu_0_jtag_debug_module_writedata;
  reg              d1_cpu_0_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module;
  wire    [ 24: 0] shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master;
  wire             wait_for_cpu_0_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_0_jtag_debug_module_end_xfer;
    end


  assign cpu_0_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module | cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module));
  //assign cpu_0_jtag_debug_module_readdata_from_sa = cpu_0_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_0_jtag_debug_module_readdata_from_sa = cpu_0_jtag_debug_module_readdata;

  assign cpu_0_data_master_requests_cpu_0_jtag_debug_module = ({cpu_0_data_master_address_to_slave[24 : 11] , 11'b0} == 25'h1902800) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //cpu_0_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_0_jtag_debug_module_arb_share_set_values = 1;

  //cpu_0_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_0_jtag_debug_module_non_bursting_master_requests = cpu_0_data_master_requests_cpu_0_jtag_debug_module |
    cpu_0_instruction_master_requests_cpu_0_jtag_debug_module |
    cpu_0_data_master_requests_cpu_0_jtag_debug_module |
    cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;

  //cpu_0_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_0_jtag_debug_module_any_bursting_master_saved_grant = 0;

  //cpu_0_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_0_jtag_debug_module_arb_share_counter_next_value = cpu_0_jtag_debug_module_firsttransfer ? (cpu_0_jtag_debug_module_arb_share_set_values - 1) : |cpu_0_jtag_debug_module_arb_share_counter ? (cpu_0_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_0_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_0_jtag_debug_module_allgrants = (|cpu_0_jtag_debug_module_grant_vector) |
    (|cpu_0_jtag_debug_module_grant_vector) |
    (|cpu_0_jtag_debug_module_grant_vector) |
    (|cpu_0_jtag_debug_module_grant_vector);

  //cpu_0_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_0_jtag_debug_module_end_xfer = ~(cpu_0_jtag_debug_module_waits_for_read | cpu_0_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module = cpu_0_jtag_debug_module_end_xfer & (~cpu_0_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_0_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_0_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module & cpu_0_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module & ~cpu_0_jtag_debug_module_non_bursting_master_requests);

  //cpu_0_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_0_jtag_debug_module_arb_counter_enable)
          cpu_0_jtag_debug_module_arb_share_counter <= cpu_0_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_0_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_0_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module & ~cpu_0_jtag_debug_module_non_bursting_master_requests))
          cpu_0_jtag_debug_module_slavearbiterlockenable <= |cpu_0_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_0/data_master cpu_0/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = cpu_0_jtag_debug_module_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //cpu_0_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_0_jtag_debug_module_slavearbiterlockenable2 = |cpu_0_jtag_debug_module_arb_share_counter_next_value;

  //cpu_0/data_master cpu_0/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = cpu_0_jtag_debug_module_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master cpu_0/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = cpu_0_jtag_debug_module_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master cpu_0/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = cpu_0_jtag_debug_module_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted cpu_0/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module <= cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module ? 1 : (cpu_0_jtag_debug_module_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_cpu_0_jtag_debug_module) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module & cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;

  //cpu_0_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_0_jtag_debug_module_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest;

  assign cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module = cpu_0_data_master_requests_cpu_0_jtag_debug_module & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_instruction_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module, which is an e_mux
  assign cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module = cpu_0_data_master_granted_cpu_0_jtag_debug_module & cpu_0_data_master_read & ~cpu_0_jtag_debug_module_waits_for_read;

  //cpu_0_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_0_jtag_debug_module_writedata = cpu_0_data_master_writedata;

  assign cpu_0_instruction_master_requests_cpu_0_jtag_debug_module = (({cpu_0_instruction_master_address_to_slave[24 : 11] , 11'b0} == 25'h1902800) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted cpu_0/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module <= cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module ? 1 : (cpu_0_jtag_debug_module_arbitration_holdoff_internal | ~cpu_0_data_master_requests_cpu_0_jtag_debug_module) ? 0 : last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module & cpu_0_data_master_requests_cpu_0_jtag_debug_module;

  assign cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module = cpu_0_instruction_master_requests_cpu_0_jtag_debug_module & ~((cpu_0_instruction_master_read & ((cpu_0_instruction_master_latency_counter != 0))) | cpu_0_data_master_arbiterlock);
  //local readdatavalid cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module = cpu_0_instruction_master_granted_cpu_0_jtag_debug_module & cpu_0_instruction_master_read & ~cpu_0_jtag_debug_module_waits_for_read;

  //allow new arb cycle for cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_jtag_debug_module_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock;

  //cpu_0/instruction_master assignment into master qualified-requests vector for cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_jtag_debug_module_master_qreq_vector[0] = cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;

  //cpu_0/instruction_master grant cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_instruction_master_granted_cpu_0_jtag_debug_module = cpu_0_jtag_debug_module_grant_vector[0];

  //cpu_0/instruction_master saved-grant cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module = cpu_0_jtag_debug_module_arb_winner[0] && cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;

  //cpu_0/data_master assignment into master qualified-requests vector for cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_jtag_debug_module_master_qreq_vector[1] = cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;

  //cpu_0/data_master grant cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_data_master_granted_cpu_0_jtag_debug_module = cpu_0_jtag_debug_module_grant_vector[1];

  //cpu_0/data_master saved-grant cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module = cpu_0_jtag_debug_module_arb_winner[1] && cpu_0_data_master_requests_cpu_0_jtag_debug_module;

  //cpu_0/jtag_debug_module chosen-master double-vector, which is an e_assign
  assign cpu_0_jtag_debug_module_chosen_master_double_vector = {cpu_0_jtag_debug_module_master_qreq_vector, cpu_0_jtag_debug_module_master_qreq_vector} & ({~cpu_0_jtag_debug_module_master_qreq_vector, ~cpu_0_jtag_debug_module_master_qreq_vector} + cpu_0_jtag_debug_module_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_0_jtag_debug_module_arb_winner = (cpu_0_jtag_debug_module_allow_new_arb_cycle & | cpu_0_jtag_debug_module_grant_vector) ? cpu_0_jtag_debug_module_grant_vector : cpu_0_jtag_debug_module_saved_chosen_master_vector;

  //saved cpu_0_jtag_debug_module_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_jtag_debug_module_saved_chosen_master_vector <= 0;
      else if (cpu_0_jtag_debug_module_allow_new_arb_cycle)
          cpu_0_jtag_debug_module_saved_chosen_master_vector <= |cpu_0_jtag_debug_module_grant_vector ? cpu_0_jtag_debug_module_grant_vector : cpu_0_jtag_debug_module_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_0_jtag_debug_module_grant_vector = {(cpu_0_jtag_debug_module_chosen_master_double_vector[1] | cpu_0_jtag_debug_module_chosen_master_double_vector[3]),
    (cpu_0_jtag_debug_module_chosen_master_double_vector[0] | cpu_0_jtag_debug_module_chosen_master_double_vector[2])};

  //cpu_0/jtag_debug_module chosen master rotated left, which is an e_assign
  assign cpu_0_jtag_debug_module_chosen_master_rot_left = (cpu_0_jtag_debug_module_arb_winner << 1) ? (cpu_0_jtag_debug_module_arb_winner << 1) : 1;

  //cpu_0/jtag_debug_module's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_jtag_debug_module_arb_addend <= 1;
      else if (|cpu_0_jtag_debug_module_grant_vector)
          cpu_0_jtag_debug_module_arb_addend <= cpu_0_jtag_debug_module_end_xfer? cpu_0_jtag_debug_module_chosen_master_rot_left : cpu_0_jtag_debug_module_grant_vector;
    end


  assign cpu_0_jtag_debug_module_begintransfer = cpu_0_jtag_debug_module_begins_xfer;
  //assign cpu_0_jtag_debug_module_resetrequest_from_sa = cpu_0_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_0_jtag_debug_module_resetrequest_from_sa = cpu_0_jtag_debug_module_resetrequest;

  assign cpu_0_jtag_debug_module_chipselect = cpu_0_data_master_granted_cpu_0_jtag_debug_module | cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  //cpu_0_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_0_jtag_debug_module_firsttransfer = cpu_0_jtag_debug_module_begins_xfer ? cpu_0_jtag_debug_module_unreg_firsttransfer : cpu_0_jtag_debug_module_reg_firsttransfer;

  //cpu_0_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_0_jtag_debug_module_unreg_firsttransfer = ~(cpu_0_jtag_debug_module_slavearbiterlockenable & cpu_0_jtag_debug_module_any_continuerequest);

  //cpu_0_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_0_jtag_debug_module_begins_xfer)
          cpu_0_jtag_debug_module_reg_firsttransfer <= cpu_0_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_0_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_0_jtag_debug_module_beginbursttransfer_internal = cpu_0_jtag_debug_module_begins_xfer;

  //cpu_0_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_0_jtag_debug_module_arbitration_holdoff_internal = cpu_0_jtag_debug_module_begins_xfer & cpu_0_jtag_debug_module_firsttransfer;

  //cpu_0_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_0_jtag_debug_module_write = cpu_0_data_master_granted_cpu_0_jtag_debug_module & cpu_0_data_master_write;

  assign shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //cpu_0_jtag_debug_module_address mux, which is an e_mux
  assign cpu_0_jtag_debug_module_address = (cpu_0_data_master_granted_cpu_0_jtag_debug_module)? (shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master >> 2) :
    (shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master >> 2);

  assign shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master = cpu_0_instruction_master_address_to_slave;
  //d1_cpu_0_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_0_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_0_jtag_debug_module_end_xfer <= cpu_0_jtag_debug_module_end_xfer;
    end


  //cpu_0_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_0_jtag_debug_module_waits_for_read = cpu_0_jtag_debug_module_in_a_read_cycle & cpu_0_jtag_debug_module_begins_xfer;

  //cpu_0_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_0_jtag_debug_module_in_a_read_cycle = (cpu_0_data_master_granted_cpu_0_jtag_debug_module & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_cpu_0_jtag_debug_module & cpu_0_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_0_jtag_debug_module_in_a_read_cycle;

  //cpu_0_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_0_jtag_debug_module_waits_for_write = cpu_0_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_0_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_0_jtag_debug_module_in_a_write_cycle = cpu_0_data_master_granted_cpu_0_jtag_debug_module & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_0_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_0_jtag_debug_module_counter = 0;
  //cpu_0_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_0_jtag_debug_module_byteenable = (cpu_0_data_master_granted_cpu_0_jtag_debug_module)? cpu_0_data_master_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_0_jtag_debug_module_debugaccess = (cpu_0_data_master_granted_cpu_0_jtag_debug_module)? cpu_0_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_0/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_cpu_0_jtag_debug_module + cpu_0_instruction_master_granted_cpu_0_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module + cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_0_custom_instruction_master_arbitrator (
                                                    // inputs:
                                                     clk,
                                                     cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa,
                                                     cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa,
                                                     cpu_0_custom_instruction_master_multi_start,
                                                     reset_n,

                                                    // outputs:
                                                     cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select,
                                                     cpu_0_custom_instruction_master_multi_done,
                                                     cpu_0_custom_instruction_master_multi_result,
                                                     cpu_0_custom_instruction_master_reset_n,
                                                     cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1
                                                  )
;

  output           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select;
  output           cpu_0_custom_instruction_master_multi_done;
  output  [ 31: 0] cpu_0_custom_instruction_master_multi_result;
  output           cpu_0_custom_instruction_master_reset_n;
  output           cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1;
  input            clk;
  input            cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  input   [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  input            cpu_0_custom_instruction_master_multi_start;
  input            reset_n;

  wire             cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select;
  wire             cpu_0_custom_instruction_master_multi_done;
  wire    [ 31: 0] cpu_0_custom_instruction_master_multi_result;
  wire             cpu_0_custom_instruction_master_reset_n;
  wire             cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1;
  assign cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select = 1'b1;
  assign cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1 = cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select & cpu_0_custom_instruction_master_multi_start;
  //cpu_0_custom_instruction_master_multi_result mux, which is an e_mux
  assign cpu_0_custom_instruction_master_multi_result = {32 {cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select}} & cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;

  //multi_done mux, which is an e_mux
  assign cpu_0_custom_instruction_master_multi_done = {1 {cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select}} & cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;

  //cpu_0_custom_instruction_master_reset_n local reset_n, which is an e_assign
  assign cpu_0_custom_instruction_master_reset_n = reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_0_data_master_arbitrator (
                                      // inputs:
                                       clk,
                                       cpu_0_data_master_address,
                                       cpu_0_data_master_byteenable,
                                       cpu_0_data_master_byteenable_nios_system_clock_3_in,
                                       cpu_0_data_master_byteenable_nios_system_clock_9_in,
                                       cpu_0_data_master_byteenable_sram_0_avalon_sram_slave,
                                       cpu_0_data_master_granted_cpu_0_jtag_debug_module,
                                       cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave,
                                       cpu_0_data_master_granted_keys_s1,
                                       cpu_0_data_master_granted_mailbox_0_s1,
                                       cpu_0_data_master_granted_mailbox_1_s1,
                                       cpu_0_data_master_granted_mailbox_2_s1,
                                       cpu_0_data_master_granted_mailbox_3_s1,
                                       cpu_0_data_master_granted_nios_system_clock_3_in,
                                       cpu_0_data_master_granted_nios_system_clock_9_in,
                                       cpu_0_data_master_granted_onchip_memory2_0_s1,
                                       cpu_0_data_master_granted_onchip_memory2_1_s1,
                                       cpu_0_data_master_granted_onchip_memory2_2_s1,
                                       cpu_0_data_master_granted_onchip_memory2_3_s1,
                                       cpu_0_data_master_granted_performance_counter_0_control_slave,
                                       cpu_0_data_master_granted_sram_0_avalon_sram_slave,
                                       cpu_0_data_master_granted_sysid_control_slave,
                                       cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module,
                                       cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave,
                                       cpu_0_data_master_qualified_request_keys_s1,
                                       cpu_0_data_master_qualified_request_mailbox_0_s1,
                                       cpu_0_data_master_qualified_request_mailbox_1_s1,
                                       cpu_0_data_master_qualified_request_mailbox_2_s1,
                                       cpu_0_data_master_qualified_request_mailbox_3_s1,
                                       cpu_0_data_master_qualified_request_nios_system_clock_3_in,
                                       cpu_0_data_master_qualified_request_nios_system_clock_9_in,
                                       cpu_0_data_master_qualified_request_onchip_memory2_0_s1,
                                       cpu_0_data_master_qualified_request_onchip_memory2_1_s1,
                                       cpu_0_data_master_qualified_request_onchip_memory2_2_s1,
                                       cpu_0_data_master_qualified_request_onchip_memory2_3_s1,
                                       cpu_0_data_master_qualified_request_performance_counter_0_control_slave,
                                       cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave,
                                       cpu_0_data_master_qualified_request_sysid_control_slave,
                                       cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_0_data_master_read,
                                       cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module,
                                       cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave,
                                       cpu_0_data_master_read_data_valid_keys_s1,
                                       cpu_0_data_master_read_data_valid_mailbox_0_s1,
                                       cpu_0_data_master_read_data_valid_mailbox_1_s1,
                                       cpu_0_data_master_read_data_valid_mailbox_2_s1,
                                       cpu_0_data_master_read_data_valid_mailbox_3_s1,
                                       cpu_0_data_master_read_data_valid_nios_system_clock_3_in,
                                       cpu_0_data_master_read_data_valid_nios_system_clock_9_in,
                                       cpu_0_data_master_read_data_valid_onchip_memory2_0_s1,
                                       cpu_0_data_master_read_data_valid_onchip_memory2_1_s1,
                                       cpu_0_data_master_read_data_valid_onchip_memory2_2_s1,
                                       cpu_0_data_master_read_data_valid_onchip_memory2_3_s1,
                                       cpu_0_data_master_read_data_valid_performance_counter_0_control_slave,
                                       cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave,
                                       cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                       cpu_0_data_master_read_data_valid_sysid_control_slave,
                                       cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_0_data_master_requests_cpu_0_jtag_debug_module,
                                       cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave,
                                       cpu_0_data_master_requests_keys_s1,
                                       cpu_0_data_master_requests_mailbox_0_s1,
                                       cpu_0_data_master_requests_mailbox_1_s1,
                                       cpu_0_data_master_requests_mailbox_2_s1,
                                       cpu_0_data_master_requests_mailbox_3_s1,
                                       cpu_0_data_master_requests_nios_system_clock_3_in,
                                       cpu_0_data_master_requests_nios_system_clock_9_in,
                                       cpu_0_data_master_requests_onchip_memory2_0_s1,
                                       cpu_0_data_master_requests_onchip_memory2_1_s1,
                                       cpu_0_data_master_requests_onchip_memory2_2_s1,
                                       cpu_0_data_master_requests_onchip_memory2_3_s1,
                                       cpu_0_data_master_requests_performance_counter_0_control_slave,
                                       cpu_0_data_master_requests_sram_0_avalon_sram_slave,
                                       cpu_0_data_master_requests_sysid_control_slave,
                                       cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_0_data_master_write,
                                       cpu_0_data_master_writedata,
                                       cpu_0_jtag_debug_module_readdata_from_sa,
                                       d1_cpu_0_jtag_debug_module_end_xfer,
                                       d1_jtag_uart_0_avalon_jtag_slave_end_xfer,
                                       d1_keys_s1_end_xfer,
                                       d1_mailbox_0_s1_end_xfer,
                                       d1_mailbox_1_s1_end_xfer,
                                       d1_mailbox_2_s1_end_xfer,
                                       d1_mailbox_3_s1_end_xfer,
                                       d1_nios_system_clock_3_in_end_xfer,
                                       d1_nios_system_clock_9_in_end_xfer,
                                       d1_onchip_memory2_0_s1_end_xfer,
                                       d1_onchip_memory2_1_s1_end_xfer,
                                       d1_onchip_memory2_2_s1_end_xfer,
                                       d1_onchip_memory2_3_s1_end_xfer,
                                       d1_performance_counter_0_control_slave_end_xfer,
                                       d1_sram_0_avalon_sram_slave_end_xfer,
                                       d1_sysid_control_slave_end_xfer,
                                       d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer,
                                       jtag_uart_0_avalon_jtag_slave_irq_from_sa,
                                       jtag_uart_0_avalon_jtag_slave_readdata_from_sa,
                                       jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa,
                                       keys_s1_readdata_from_sa,
                                       mailbox_0_s1_readdata_from_sa,
                                       mailbox_1_s1_readdata_from_sa,
                                       mailbox_2_s1_readdata_from_sa,
                                       mailbox_3_s1_readdata_from_sa,
                                       nios_system_clock_3_in_readdata_from_sa,
                                       nios_system_clock_3_in_waitrequest_from_sa,
                                       nios_system_clock_9_in_readdata_from_sa,
                                       nios_system_clock_9_in_waitrequest_from_sa,
                                       onchip_memory2_0_s1_readdata_from_sa,
                                       onchip_memory2_1_s1_readdata_from_sa,
                                       onchip_memory2_2_s1_readdata_from_sa,
                                       onchip_memory2_3_s1_readdata_from_sa,
                                       performance_counter_0_control_slave_readdata_from_sa,
                                       reset_n,
                                       sram_0_avalon_sram_slave_readdata_from_sa,
                                       sysid_control_slave_readdata_from_sa,
                                       video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa,

                                      // outputs:
                                       cpu_0_data_master_address_to_slave,
                                       cpu_0_data_master_dbs_address,
                                       cpu_0_data_master_dbs_write_16,
                                       cpu_0_data_master_dbs_write_8,
                                       cpu_0_data_master_irq,
                                       cpu_0_data_master_latency_counter,
                                       cpu_0_data_master_readdata,
                                       cpu_0_data_master_readdatavalid,
                                       cpu_0_data_master_waitrequest
                                    )
;

  output  [ 24: 0] cpu_0_data_master_address_to_slave;
  output  [  1: 0] cpu_0_data_master_dbs_address;
  output  [ 15: 0] cpu_0_data_master_dbs_write_16;
  output  [  7: 0] cpu_0_data_master_dbs_write_8;
  output  [ 31: 0] cpu_0_data_master_irq;
  output           cpu_0_data_master_latency_counter;
  output  [ 31: 0] cpu_0_data_master_readdata;
  output           cpu_0_data_master_readdatavalid;
  output           cpu_0_data_master_waitrequest;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input   [  1: 0] cpu_0_data_master_byteenable_nios_system_clock_3_in;
  input            cpu_0_data_master_byteenable_nios_system_clock_9_in;
  input   [  1: 0] cpu_0_data_master_byteenable_sram_0_avalon_sram_slave;
  input            cpu_0_data_master_granted_cpu_0_jtag_debug_module;
  input            cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave;
  input            cpu_0_data_master_granted_keys_s1;
  input            cpu_0_data_master_granted_mailbox_0_s1;
  input            cpu_0_data_master_granted_mailbox_1_s1;
  input            cpu_0_data_master_granted_mailbox_2_s1;
  input            cpu_0_data_master_granted_mailbox_3_s1;
  input            cpu_0_data_master_granted_nios_system_clock_3_in;
  input            cpu_0_data_master_granted_nios_system_clock_9_in;
  input            cpu_0_data_master_granted_onchip_memory2_0_s1;
  input            cpu_0_data_master_granted_onchip_memory2_1_s1;
  input            cpu_0_data_master_granted_onchip_memory2_2_s1;
  input            cpu_0_data_master_granted_onchip_memory2_3_s1;
  input            cpu_0_data_master_granted_performance_counter_0_control_slave;
  input            cpu_0_data_master_granted_sram_0_avalon_sram_slave;
  input            cpu_0_data_master_granted_sysid_control_slave;
  input            cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  input            cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave;
  input            cpu_0_data_master_qualified_request_keys_s1;
  input            cpu_0_data_master_qualified_request_mailbox_0_s1;
  input            cpu_0_data_master_qualified_request_mailbox_1_s1;
  input            cpu_0_data_master_qualified_request_mailbox_2_s1;
  input            cpu_0_data_master_qualified_request_mailbox_3_s1;
  input            cpu_0_data_master_qualified_request_nios_system_clock_3_in;
  input            cpu_0_data_master_qualified_request_nios_system_clock_9_in;
  input            cpu_0_data_master_qualified_request_onchip_memory2_0_s1;
  input            cpu_0_data_master_qualified_request_onchip_memory2_1_s1;
  input            cpu_0_data_master_qualified_request_onchip_memory2_2_s1;
  input            cpu_0_data_master_qualified_request_onchip_memory2_3_s1;
  input            cpu_0_data_master_qualified_request_performance_counter_0_control_slave;
  input            cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave;
  input            cpu_0_data_master_qualified_request_sysid_control_slave;
  input            cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module;
  input            cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  input            cpu_0_data_master_read_data_valid_keys_s1;
  input            cpu_0_data_master_read_data_valid_mailbox_0_s1;
  input            cpu_0_data_master_read_data_valid_mailbox_1_s1;
  input            cpu_0_data_master_read_data_valid_mailbox_2_s1;
  input            cpu_0_data_master_read_data_valid_mailbox_3_s1;
  input            cpu_0_data_master_read_data_valid_nios_system_clock_3_in;
  input            cpu_0_data_master_read_data_valid_nios_system_clock_9_in;
  input            cpu_0_data_master_read_data_valid_onchip_memory2_0_s1;
  input            cpu_0_data_master_read_data_valid_onchip_memory2_1_s1;
  input            cpu_0_data_master_read_data_valid_onchip_memory2_2_s1;
  input            cpu_0_data_master_read_data_valid_onchip_memory2_3_s1;
  input            cpu_0_data_master_read_data_valid_performance_counter_0_control_slave;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_read_data_valid_sysid_control_slave;
  input            cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  input            cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;
  input            cpu_0_data_master_requests_keys_s1;
  input            cpu_0_data_master_requests_mailbox_0_s1;
  input            cpu_0_data_master_requests_mailbox_1_s1;
  input            cpu_0_data_master_requests_mailbox_2_s1;
  input            cpu_0_data_master_requests_mailbox_3_s1;
  input            cpu_0_data_master_requests_nios_system_clock_3_in;
  input            cpu_0_data_master_requests_nios_system_clock_9_in;
  input            cpu_0_data_master_requests_onchip_memory2_0_s1;
  input            cpu_0_data_master_requests_onchip_memory2_1_s1;
  input            cpu_0_data_master_requests_onchip_memory2_2_s1;
  input            cpu_0_data_master_requests_onchip_memory2_3_s1;
  input            cpu_0_data_master_requests_performance_counter_0_control_slave;
  input            cpu_0_data_master_requests_sram_0_avalon_sram_slave;
  input            cpu_0_data_master_requests_sysid_control_slave;
  input            cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 31: 0] cpu_0_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_0_jtag_debug_module_end_xfer;
  input            d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  input            d1_keys_s1_end_xfer;
  input            d1_mailbox_0_s1_end_xfer;
  input            d1_mailbox_1_s1_end_xfer;
  input            d1_mailbox_2_s1_end_xfer;
  input            d1_mailbox_3_s1_end_xfer;
  input            d1_nios_system_clock_3_in_end_xfer;
  input            d1_nios_system_clock_9_in_end_xfer;
  input            d1_onchip_memory2_0_s1_end_xfer;
  input            d1_onchip_memory2_1_s1_end_xfer;
  input            d1_onchip_memory2_2_s1_end_xfer;
  input            d1_onchip_memory2_3_s1_end_xfer;
  input            d1_performance_counter_0_control_slave_end_xfer;
  input            d1_sram_0_avalon_sram_slave_end_xfer;
  input            d1_sysid_control_slave_end_xfer;
  input            d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer;
  input            jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  input   [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  input   [ 31: 0] keys_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_0_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_1_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_2_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_3_s1_readdata_from_sa;
  input   [ 15: 0] nios_system_clock_3_in_readdata_from_sa;
  input            nios_system_clock_3_in_waitrequest_from_sa;
  input   [  7: 0] nios_system_clock_9_in_readdata_from_sa;
  input            nios_system_clock_9_in_waitrequest_from_sa;
  input   [ 31: 0] onchip_memory2_0_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_1_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_2_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_3_s1_readdata_from_sa;
  input   [ 31: 0] performance_counter_0_control_slave_readdata_from_sa;
  input            reset_n;
  input   [ 15: 0] sram_0_avalon_sram_slave_readdata_from_sa;
  input   [ 31: 0] sysid_control_slave_readdata_from_sa;
  input   [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] cpu_0_data_master_address_last_time;
  wire    [ 24: 0] cpu_0_data_master_address_to_slave;
  reg     [  3: 0] cpu_0_data_master_byteenable_last_time;
  reg     [  1: 0] cpu_0_data_master_dbs_address;
  wire    [  1: 0] cpu_0_data_master_dbs_increment;
  reg     [  1: 0] cpu_0_data_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_0_data_master_dbs_rdv_counter_inc;
  wire    [ 15: 0] cpu_0_data_master_dbs_write_16;
  wire    [  7: 0] cpu_0_data_master_dbs_write_8;
  wire    [ 31: 0] cpu_0_data_master_irq;
  wire             cpu_0_data_master_is_granted_some_slave;
  reg              cpu_0_data_master_latency_counter;
  wire    [  1: 0] cpu_0_data_master_next_dbs_rdv_counter;
  reg              cpu_0_data_master_read_but_no_slave_selected;
  reg              cpu_0_data_master_read_last_time;
  wire    [ 31: 0] cpu_0_data_master_readdata;
  wire             cpu_0_data_master_readdatavalid;
  wire             cpu_0_data_master_run;
  wire             cpu_0_data_master_waitrequest;
  reg              cpu_0_data_master_write_last_time;
  reg     [ 31: 0] cpu_0_data_master_writedata_last_time;
  reg     [ 15: 0] dbs_16_reg_segment_0;
  reg     [  7: 0] dbs_8_reg_segment_0;
  reg     [  7: 0] dbs_8_reg_segment_1;
  reg     [  7: 0] dbs_8_reg_segment_2;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire             p1_cpu_0_data_master_latency_counter;
  wire    [ 15: 0] p1_dbs_16_reg_segment_0;
  wire    [  7: 0] p1_dbs_8_reg_segment_0;
  wire    [  7: 0] p1_dbs_8_reg_segment_1;
  wire    [  7: 0] p1_dbs_8_reg_segment_2;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_0_data_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  wire             r_3;
  wire             r_4;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module | ~cpu_0_data_master_requests_cpu_0_jtag_debug_module) & (cpu_0_data_master_granted_cpu_0_jtag_debug_module | ~cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module) & ((~cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module | ~cpu_0_data_master_read | (1 & ~d1_cpu_0_jtag_debug_module_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave | ~cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave) & ((~cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & ~jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa & (cpu_0_data_master_read | cpu_0_data_master_write)))) & ((~cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & ~jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa & (cpu_0_data_master_read | cpu_0_data_master_write)))) & 1 & (cpu_0_data_master_qualified_request_keys_s1 | ~cpu_0_data_master_requests_keys_s1) & (cpu_0_data_master_granted_keys_s1 | ~cpu_0_data_master_qualified_request_keys_s1) & ((~cpu_0_data_master_qualified_request_keys_s1 | ~cpu_0_data_master_read | (1 & ~d1_keys_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_keys_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_mailbox_0_s1 | ~cpu_0_data_master_requests_mailbox_0_s1) & (cpu_0_data_master_granted_mailbox_0_s1 | ~cpu_0_data_master_qualified_request_mailbox_0_s1) & ((~cpu_0_data_master_qualified_request_mailbox_0_s1 | ~cpu_0_data_master_read | (1 & ~d1_mailbox_0_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_mailbox_0_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1;

  //cascaded wait assignment, which is an e_assign
  assign cpu_0_data_master_run = r_0 & r_1 & r_2 & r_3 & r_4;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = (cpu_0_data_master_qualified_request_mailbox_1_s1 | ~cpu_0_data_master_requests_mailbox_1_s1) & (cpu_0_data_master_granted_mailbox_1_s1 | ~cpu_0_data_master_qualified_request_mailbox_1_s1) & ((~cpu_0_data_master_qualified_request_mailbox_1_s1 | ~cpu_0_data_master_read | (1 & ~d1_mailbox_1_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_mailbox_1_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_mailbox_2_s1 | ~cpu_0_data_master_requests_mailbox_2_s1) & (cpu_0_data_master_granted_mailbox_2_s1 | ~cpu_0_data_master_qualified_request_mailbox_2_s1) & ((~cpu_0_data_master_qualified_request_mailbox_2_s1 | ~cpu_0_data_master_read | (1 & ~d1_mailbox_2_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_mailbox_2_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_mailbox_3_s1 | ~cpu_0_data_master_requests_mailbox_3_s1) & (cpu_0_data_master_granted_mailbox_3_s1 | ~cpu_0_data_master_qualified_request_mailbox_3_s1) & ((~cpu_0_data_master_qualified_request_mailbox_3_s1 | ~cpu_0_data_master_read | (1 & ~d1_mailbox_3_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_mailbox_3_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_nios_system_clock_3_in | (cpu_0_data_master_write & !cpu_0_data_master_byteenable_nios_system_clock_3_in & cpu_0_data_master_dbs_address[1]) | ~cpu_0_data_master_requests_nios_system_clock_3_in) & ((~cpu_0_data_master_qualified_request_nios_system_clock_3_in | ~cpu_0_data_master_read | (1 & ~nios_system_clock_3_in_waitrequest_from_sa & (cpu_0_data_master_dbs_address[1]) & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_nios_system_clock_3_in | ~cpu_0_data_master_write | (1 & ~nios_system_clock_3_in_waitrequest_from_sa & (cpu_0_data_master_dbs_address[1]) & cpu_0_data_master_write)));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & ((cpu_0_data_master_qualified_request_nios_system_clock_9_in | ((cpu_0_data_master_write & !cpu_0_data_master_byteenable_nios_system_clock_9_in & cpu_0_data_master_dbs_address[1] & cpu_0_data_master_dbs_address[0])) | ~cpu_0_data_master_requests_nios_system_clock_9_in)) & ((~cpu_0_data_master_qualified_request_nios_system_clock_9_in | ~cpu_0_data_master_read | (1 & ~nios_system_clock_9_in_waitrequest_from_sa & (cpu_0_data_master_dbs_address[1] & cpu_0_data_master_dbs_address[0]) & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_nios_system_clock_9_in | ~cpu_0_data_master_write | (1 & ~nios_system_clock_9_in_waitrequest_from_sa & (cpu_0_data_master_dbs_address[1] & cpu_0_data_master_dbs_address[0]) & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_onchip_memory2_0_s1 | ~cpu_0_data_master_requests_onchip_memory2_0_s1) & (cpu_0_data_master_granted_onchip_memory2_0_s1 | ~cpu_0_data_master_qualified_request_onchip_memory2_0_s1) & ((~cpu_0_data_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write)))) & ((~cpu_0_data_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write)))) & 1 & (cpu_0_data_master_qualified_request_onchip_memory2_1_s1 | ~cpu_0_data_master_requests_onchip_memory2_1_s1) & (cpu_0_data_master_granted_onchip_memory2_1_s1 | ~cpu_0_data_master_qualified_request_onchip_memory2_1_s1) & ((~cpu_0_data_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write)))) & ((~cpu_0_data_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write)))) & 1 & (cpu_0_data_master_qualified_request_onchip_memory2_2_s1 | ~cpu_0_data_master_requests_onchip_memory2_2_s1) & (cpu_0_data_master_granted_onchip_memory2_2_s1 | ~cpu_0_data_master_qualified_request_onchip_memory2_2_s1) & ((~cpu_0_data_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write)))) & ((~cpu_0_data_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write)))) & 1;

  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = (cpu_0_data_master_qualified_request_onchip_memory2_3_s1 | ~cpu_0_data_master_requests_onchip_memory2_3_s1) & (cpu_0_data_master_granted_onchip_memory2_3_s1 | ~cpu_0_data_master_qualified_request_onchip_memory2_3_s1) & ((~cpu_0_data_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write)))) & ((~cpu_0_data_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write)))) & 1 & (cpu_0_data_master_qualified_request_performance_counter_0_control_slave | ~cpu_0_data_master_requests_performance_counter_0_control_slave) & (cpu_0_data_master_granted_performance_counter_0_control_slave | ~cpu_0_data_master_qualified_request_performance_counter_0_control_slave) & ((~cpu_0_data_master_qualified_request_performance_counter_0_control_slave | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write)))) & ((~cpu_0_data_master_qualified_request_performance_counter_0_control_slave | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write)))) & 1 & (cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave | (cpu_0_data_master_write & !cpu_0_data_master_byteenable_sram_0_avalon_sram_slave & cpu_0_data_master_dbs_address[1]) | ~cpu_0_data_master_requests_sram_0_avalon_sram_slave) & (cpu_0_data_master_granted_sram_0_avalon_sram_slave | ~cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave) & ((~cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_0_data_master_read | (1 & (cpu_0_data_master_dbs_address[1]) & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_0_data_master_write | (1 & (cpu_0_data_master_dbs_address[1]) & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_sysid_control_slave | ~cpu_0_data_master_requests_sysid_control_slave) & (cpu_0_data_master_granted_sysid_control_slave | ~cpu_0_data_master_qualified_request_sysid_control_slave) & ((~cpu_0_data_master_qualified_request_sysid_control_slave | ~cpu_0_data_master_read | (1 & ~d1_sysid_control_slave_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_sysid_control_slave | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write)));

  //r_4 master_run cascaded wait assignment, which is an e_assign
  assign r_4 = 1 & (cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) & (cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave | ~cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave) & ((~cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write)))) & ((~cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & (cpu_0_data_master_read | cpu_0_data_master_write))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_0_data_master_address_to_slave = cpu_0_data_master_address[24 : 0];

  //cpu_0_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_read_but_no_slave_selected <= 0;
      else 
        cpu_0_data_master_read_but_no_slave_selected <= cpu_0_data_master_read & cpu_0_data_master_run & ~cpu_0_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_0_data_master_is_granted_some_slave = cpu_0_data_master_granted_cpu_0_jtag_debug_module |
    cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave |
    cpu_0_data_master_granted_keys_s1 |
    cpu_0_data_master_granted_mailbox_0_s1 |
    cpu_0_data_master_granted_mailbox_1_s1 |
    cpu_0_data_master_granted_mailbox_2_s1 |
    cpu_0_data_master_granted_mailbox_3_s1 |
    cpu_0_data_master_granted_nios_system_clock_3_in |
    cpu_0_data_master_granted_nios_system_clock_9_in |
    cpu_0_data_master_granted_onchip_memory2_0_s1 |
    cpu_0_data_master_granted_onchip_memory2_1_s1 |
    cpu_0_data_master_granted_onchip_memory2_2_s1 |
    cpu_0_data_master_granted_onchip_memory2_3_s1 |
    cpu_0_data_master_granted_performance_counter_0_control_slave |
    cpu_0_data_master_granted_sram_0_avalon_sram_slave |
    cpu_0_data_master_granted_sysid_control_slave |
    cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_0_data_master_readdatavalid = cpu_0_data_master_read_data_valid_onchip_memory2_0_s1 |
    cpu_0_data_master_read_data_valid_onchip_memory2_1_s1 |
    cpu_0_data_master_read_data_valid_onchip_memory2_2_s1 |
    cpu_0_data_master_read_data_valid_onchip_memory2_3_s1 |
    cpu_0_data_master_read_data_valid_performance_counter_0_control_slave |
    (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave & dbs_rdv_counter_overflow) |
    cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_0_data_master_readdatavalid = cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_keys_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_mailbox_0_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_mailbox_1_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_mailbox_2_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_mailbox_3_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    (cpu_0_data_master_read_data_valid_nios_system_clock_3_in & dbs_counter_overflow) |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    (cpu_0_data_master_read_data_valid_nios_system_clock_9_in & dbs_counter_overflow) |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_sysid_control_slave |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid;

  //cpu_0/data_master readdata mux, which is an e_mux
  assign cpu_0_data_master_readdata = ({32 {~(cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module & cpu_0_data_master_read)}} | cpu_0_jtag_debug_module_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_read)}} | jtag_uart_0_avalon_jtag_slave_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_keys_s1 & cpu_0_data_master_read)}} | keys_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_mailbox_0_s1 & cpu_0_data_master_read)}} | mailbox_0_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_mailbox_1_s1 & cpu_0_data_master_read)}} | mailbox_1_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_mailbox_2_s1 & cpu_0_data_master_read)}} | mailbox_2_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_mailbox_3_s1 & cpu_0_data_master_read)}} | mailbox_3_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_nios_system_clock_3_in & cpu_0_data_master_read)}} | {nios_system_clock_3_in_readdata_from_sa[15 : 0],
    dbs_16_reg_segment_0}) &
    ({32 {~(cpu_0_data_master_qualified_request_nios_system_clock_9_in & cpu_0_data_master_read)}} | {nios_system_clock_9_in_readdata_from_sa[7 : 0],
    dbs_8_reg_segment_2,
    dbs_8_reg_segment_1,
    dbs_8_reg_segment_0}) &
    ({32 {~cpu_0_data_master_read_data_valid_onchip_memory2_0_s1}} | onchip_memory2_0_s1_readdata_from_sa) &
    ({32 {~cpu_0_data_master_read_data_valid_onchip_memory2_1_s1}} | onchip_memory2_1_s1_readdata_from_sa) &
    ({32 {~cpu_0_data_master_read_data_valid_onchip_memory2_2_s1}} | onchip_memory2_2_s1_readdata_from_sa) &
    ({32 {~cpu_0_data_master_read_data_valid_onchip_memory2_3_s1}} | onchip_memory2_3_s1_readdata_from_sa) &
    ({32 {~cpu_0_data_master_read_data_valid_performance_counter_0_control_slave}} | performance_counter_0_control_slave_readdata_from_sa) &
    ({32 {~cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave}} | {sram_0_avalon_sram_slave_readdata_from_sa[15 : 0],
    dbs_latent_16_reg_segment_0}) &
    ({32 {~(cpu_0_data_master_qualified_request_sysid_control_slave & cpu_0_data_master_read)}} | sysid_control_slave_readdata_from_sa) &
    ({32 {~cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave}} | video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_0_data_master_waitrequest = ~cpu_0_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_latency_counter <= 0;
      else 
        cpu_0_data_master_latency_counter <= p1_cpu_0_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_0_data_master_latency_counter = ((cpu_0_data_master_run & cpu_0_data_master_read))? latency_load_value :
    (cpu_0_data_master_latency_counter)? cpu_0_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({1 {cpu_0_data_master_requests_onchip_memory2_0_s1}} & 1) |
    ({1 {cpu_0_data_master_requests_onchip_memory2_1_s1}} & 1) |
    ({1 {cpu_0_data_master_requests_onchip_memory2_2_s1}} & 1) |
    ({1 {cpu_0_data_master_requests_onchip_memory2_3_s1}} & 1) |
    ({1 {cpu_0_data_master_requests_performance_counter_0_control_slave}} & 1) |
    ({1 {cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave}} & 1);

  //irq assign, which is an e_assign
  assign cpu_0_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    jtag_uart_0_avalon_jtag_slave_irq_from_sa,
    1'b0};

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (((~0) & cpu_0_data_master_requests_nios_system_clock_3_in & cpu_0_data_master_write & !cpu_0_data_master_byteenable_nios_system_clock_3_in)) |
    (cpu_0_data_master_granted_nios_system_clock_3_in & cpu_0_data_master_read & 1 & 1 & ~nios_system_clock_3_in_waitrequest_from_sa) |
    (cpu_0_data_master_granted_nios_system_clock_3_in & cpu_0_data_master_write & 1 & 1 & ~nios_system_clock_3_in_waitrequest_from_sa) |
    (((~0) & cpu_0_data_master_requests_nios_system_clock_9_in & cpu_0_data_master_write & !cpu_0_data_master_byteenable_nios_system_clock_9_in)) |
    (cpu_0_data_master_granted_nios_system_clock_9_in & cpu_0_data_master_read & 1 & 1 & ~nios_system_clock_9_in_waitrequest_from_sa) |
    (cpu_0_data_master_granted_nios_system_clock_9_in & cpu_0_data_master_write & 1 & 1 & ~nios_system_clock_9_in_waitrequest_from_sa) |
    (((~0) & cpu_0_data_master_requests_sram_0_avalon_sram_slave & cpu_0_data_master_write & !cpu_0_data_master_byteenable_sram_0_avalon_sram_slave)) |
    (cpu_0_data_master_granted_sram_0_avalon_sram_slave & cpu_0_data_master_read & 1 & 1) |
    (cpu_0_data_master_granted_sram_0_avalon_sram_slave & cpu_0_data_master_write & 1 & 1);

  //input to dbs-16 stored 0, which is an e_mux
  assign p1_dbs_16_reg_segment_0 = nios_system_clock_3_in_readdata_from_sa;

  //dbs register for dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_16_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_0_data_master_dbs_address[1]) == 0))
          dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
    end


  //mux write dbs 1, which is an e_mux
  assign cpu_0_data_master_dbs_write_16 = (cpu_0_data_master_dbs_address[1])? cpu_0_data_master_writedata[31 : 16] :
    (~(cpu_0_data_master_dbs_address[1]))? cpu_0_data_master_writedata[15 : 0] :
    (cpu_0_data_master_dbs_address[1])? cpu_0_data_master_writedata[31 : 16] :
    cpu_0_data_master_writedata[15 : 0];

  //dbs count increment, which is an e_mux
  assign cpu_0_data_master_dbs_increment = (cpu_0_data_master_requests_nios_system_clock_3_in)? 2 :
    (cpu_0_data_master_requests_nios_system_clock_9_in)? 1 :
    (cpu_0_data_master_requests_sram_0_avalon_sram_slave)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_0_data_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_0_data_master_dbs_address + cpu_0_data_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_0_data_master_dbs_address <= next_dbs_address;
    end


  //input to dbs-8 stored 0, which is an e_mux
  assign p1_dbs_8_reg_segment_0 = nios_system_clock_9_in_readdata_from_sa;

  //dbs register for dbs-8 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_0_data_master_dbs_address[1 : 0]) == 0))
          dbs_8_reg_segment_0 <= p1_dbs_8_reg_segment_0;
    end


  //input to dbs-8 stored 1, which is an e_mux
  assign p1_dbs_8_reg_segment_1 = nios_system_clock_9_in_readdata_from_sa;

  //dbs register for dbs-8 segment 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_1 <= 0;
      else if (dbs_count_enable & ((cpu_0_data_master_dbs_address[1 : 0]) == 1))
          dbs_8_reg_segment_1 <= p1_dbs_8_reg_segment_1;
    end


  //input to dbs-8 stored 2, which is an e_mux
  assign p1_dbs_8_reg_segment_2 = nios_system_clock_9_in_readdata_from_sa;

  //dbs register for dbs-8 segment 2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_2 <= 0;
      else if (dbs_count_enable & ((cpu_0_data_master_dbs_address[1 : 0]) == 2))
          dbs_8_reg_segment_2 <= p1_dbs_8_reg_segment_2;
    end


  //mux write dbs 2, which is an e_mux
  assign cpu_0_data_master_dbs_write_8 = ((cpu_0_data_master_dbs_address[1 : 0] == 0))? cpu_0_data_master_writedata[7 : 0] :
    ((cpu_0_data_master_dbs_address[1 : 0] == 1))? cpu_0_data_master_writedata[15 : 8] :
    ((cpu_0_data_master_dbs_address[1 : 0] == 2))? cpu_0_data_master_writedata[23 : 16] :
    cpu_0_data_master_writedata[31 : 24];

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = sram_0_avalon_sram_slave_readdata_from_sa;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_0_data_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_0_data_master_next_dbs_rdv_counter = cpu_0_data_master_dbs_rdv_counter + cpu_0_data_master_dbs_rdv_counter_inc;

  //cpu_0_data_master_rdv_inc_mux, which is an e_mux
  assign cpu_0_data_master_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_0_data_master_dbs_rdv_counter <= cpu_0_data_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_0_data_master_dbs_rdv_counter[1] & ~cpu_0_data_master_next_dbs_rdv_counter[1];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_0_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_address_last_time <= 0;
      else 
        cpu_0_data_master_address_last_time <= cpu_0_data_master_address;
    end


  //cpu_0/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_0_data_master_waitrequest & (cpu_0_data_master_read | cpu_0_data_master_write);
    end


  //cpu_0_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_data_master_address != cpu_0_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_0_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_0_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_byteenable_last_time <= 0;
      else 
        cpu_0_data_master_byteenable_last_time <= cpu_0_data_master_byteenable;
    end


  //cpu_0_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_data_master_byteenable != cpu_0_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_0_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_0_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_read_last_time <= 0;
      else 
        cpu_0_data_master_read_last_time <= cpu_0_data_master_read;
    end


  //cpu_0_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_data_master_read != cpu_0_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_0_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_0_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_write_last_time <= 0;
      else 
        cpu_0_data_master_write_last_time <= cpu_0_data_master_write;
    end


  //cpu_0_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_data_master_write != cpu_0_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_0_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_0_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_writedata_last_time <= 0;
      else 
        cpu_0_data_master_writedata_last_time <= cpu_0_data_master_writedata;
    end


  //cpu_0_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_data_master_writedata != cpu_0_data_master_writedata_last_time) & cpu_0_data_master_write)
        begin
          $write("%0d ns: cpu_0_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_0_instruction_master_arbitrator (
                                             // inputs:
                                              clk,
                                              cpu_0_instruction_master_address,
                                              cpu_0_instruction_master_granted_cpu_0_jtag_debug_module,
                                              cpu_0_instruction_master_granted_nios_system_clock_2_in,
                                              cpu_0_instruction_master_granted_onchip_memory2_0_s1,
                                              cpu_0_instruction_master_granted_onchip_memory2_1_s1,
                                              cpu_0_instruction_master_granted_onchip_memory2_2_s1,
                                              cpu_0_instruction_master_granted_onchip_memory2_3_s1,
                                              cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module,
                                              cpu_0_instruction_master_qualified_request_nios_system_clock_2_in,
                                              cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1,
                                              cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1,
                                              cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1,
                                              cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1,
                                              cpu_0_instruction_master_read,
                                              cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module,
                                              cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in,
                                              cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1,
                                              cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1,
                                              cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1,
                                              cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1,
                                              cpu_0_instruction_master_requests_cpu_0_jtag_debug_module,
                                              cpu_0_instruction_master_requests_nios_system_clock_2_in,
                                              cpu_0_instruction_master_requests_onchip_memory2_0_s1,
                                              cpu_0_instruction_master_requests_onchip_memory2_1_s1,
                                              cpu_0_instruction_master_requests_onchip_memory2_2_s1,
                                              cpu_0_instruction_master_requests_onchip_memory2_3_s1,
                                              cpu_0_jtag_debug_module_readdata_from_sa,
                                              d1_cpu_0_jtag_debug_module_end_xfer,
                                              d1_nios_system_clock_2_in_end_xfer,
                                              d1_onchip_memory2_0_s1_end_xfer,
                                              d1_onchip_memory2_1_s1_end_xfer,
                                              d1_onchip_memory2_2_s1_end_xfer,
                                              d1_onchip_memory2_3_s1_end_xfer,
                                              nios_system_clock_2_in_readdata_from_sa,
                                              nios_system_clock_2_in_waitrequest_from_sa,
                                              onchip_memory2_0_s1_readdata_from_sa,
                                              onchip_memory2_1_s1_readdata_from_sa,
                                              onchip_memory2_2_s1_readdata_from_sa,
                                              onchip_memory2_3_s1_readdata_from_sa,
                                              reset_n,

                                             // outputs:
                                              cpu_0_instruction_master_address_to_slave,
                                              cpu_0_instruction_master_dbs_address,
                                              cpu_0_instruction_master_latency_counter,
                                              cpu_0_instruction_master_readdata,
                                              cpu_0_instruction_master_readdatavalid,
                                              cpu_0_instruction_master_waitrequest
                                           )
;

  output  [ 24: 0] cpu_0_instruction_master_address_to_slave;
  output  [  1: 0] cpu_0_instruction_master_dbs_address;
  output           cpu_0_instruction_master_latency_counter;
  output  [ 31: 0] cpu_0_instruction_master_readdata;
  output           cpu_0_instruction_master_readdatavalid;
  output           cpu_0_instruction_master_waitrequest;
  input            clk;
  input   [ 24: 0] cpu_0_instruction_master_address;
  input            cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  input            cpu_0_instruction_master_granted_nios_system_clock_2_in;
  input            cpu_0_instruction_master_granted_onchip_memory2_0_s1;
  input            cpu_0_instruction_master_granted_onchip_memory2_1_s1;
  input            cpu_0_instruction_master_granted_onchip_memory2_2_s1;
  input            cpu_0_instruction_master_granted_onchip_memory2_3_s1;
  input            cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  input            cpu_0_instruction_master_qualified_request_nios_system_clock_2_in;
  input            cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1;
  input            cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1;
  input            cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1;
  input            cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1;
  input            cpu_0_instruction_master_read;
  input            cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module;
  input            cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in;
  input            cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1;
  input            cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1;
  input            cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1;
  input            cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1;
  input            cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  input            cpu_0_instruction_master_requests_nios_system_clock_2_in;
  input            cpu_0_instruction_master_requests_onchip_memory2_0_s1;
  input            cpu_0_instruction_master_requests_onchip_memory2_1_s1;
  input            cpu_0_instruction_master_requests_onchip_memory2_2_s1;
  input            cpu_0_instruction_master_requests_onchip_memory2_3_s1;
  input   [ 31: 0] cpu_0_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_0_jtag_debug_module_end_xfer;
  input            d1_nios_system_clock_2_in_end_xfer;
  input            d1_onchip_memory2_0_s1_end_xfer;
  input            d1_onchip_memory2_1_s1_end_xfer;
  input            d1_onchip_memory2_2_s1_end_xfer;
  input            d1_onchip_memory2_3_s1_end_xfer;
  input   [ 15: 0] nios_system_clock_2_in_readdata_from_sa;
  input            nios_system_clock_2_in_waitrequest_from_sa;
  input   [ 31: 0] onchip_memory2_0_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_1_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_2_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_3_s1_readdata_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] cpu_0_instruction_master_address_last_time;
  wire    [ 24: 0] cpu_0_instruction_master_address_to_slave;
  reg     [  1: 0] cpu_0_instruction_master_dbs_address;
  wire    [  1: 0] cpu_0_instruction_master_dbs_increment;
  wire             cpu_0_instruction_master_is_granted_some_slave;
  reg              cpu_0_instruction_master_latency_counter;
  reg              cpu_0_instruction_master_read_but_no_slave_selected;
  reg              cpu_0_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_0_instruction_master_readdata;
  wire             cpu_0_instruction_master_readdatavalid;
  wire             cpu_0_instruction_master_run;
  wire             cpu_0_instruction_master_waitrequest;
  reg     [ 15: 0] dbs_16_reg_segment_0;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire             p1_cpu_0_instruction_master_latency_counter;
  wire    [ 15: 0] p1_dbs_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_0_instruction_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  wire             r_3;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module | ~cpu_0_instruction_master_requests_cpu_0_jtag_debug_module) & (cpu_0_instruction_master_granted_cpu_0_jtag_debug_module | ~cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module) & ((~cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module | ~cpu_0_instruction_master_read | (1 & ~d1_cpu_0_jtag_debug_module_end_xfer & cpu_0_instruction_master_read)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_0_instruction_master_run = r_0 & r_1 & r_2 & r_3;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_0_instruction_master_qualified_request_nios_system_clock_2_in | ~cpu_0_instruction_master_requests_nios_system_clock_2_in) & ((~cpu_0_instruction_master_qualified_request_nios_system_clock_2_in | ~cpu_0_instruction_master_read | (1 & ~nios_system_clock_2_in_waitrequest_from_sa & (cpu_0_instruction_master_dbs_address[1]) & cpu_0_instruction_master_read)));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1 | ~cpu_0_instruction_master_requests_onchip_memory2_0_s1) & (cpu_0_instruction_master_granted_onchip_memory2_0_s1 | ~cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1) & ((~cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_0_instruction_master_read) | (1 & (cpu_0_instruction_master_read)))) & 1 & (cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1 | ~cpu_0_instruction_master_requests_onchip_memory2_1_s1) & (cpu_0_instruction_master_granted_onchip_memory2_1_s1 | ~cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1) & ((~cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_0_instruction_master_read) | (1 & (cpu_0_instruction_master_read)))) & 1 & (cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1 | ~cpu_0_instruction_master_requests_onchip_memory2_2_s1) & (cpu_0_instruction_master_granted_onchip_memory2_2_s1 | ~cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1) & ((~cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_0_instruction_master_read) | (1 & (cpu_0_instruction_master_read))));

  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1 | ~cpu_0_instruction_master_requests_onchip_memory2_3_s1) & (cpu_0_instruction_master_granted_onchip_memory2_3_s1 | ~cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1) & ((~cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_0_instruction_master_read) | (1 & (cpu_0_instruction_master_read))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_0_instruction_master_address_to_slave = cpu_0_instruction_master_address[24 : 0];

  //cpu_0_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_0_instruction_master_read_but_no_slave_selected <= cpu_0_instruction_master_read & cpu_0_instruction_master_run & ~cpu_0_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_0_instruction_master_is_granted_some_slave = cpu_0_instruction_master_granted_cpu_0_jtag_debug_module |
    cpu_0_instruction_master_granted_nios_system_clock_2_in |
    cpu_0_instruction_master_granted_onchip_memory2_0_s1 |
    cpu_0_instruction_master_granted_onchip_memory2_1_s1 |
    cpu_0_instruction_master_granted_onchip_memory2_2_s1 |
    cpu_0_instruction_master_granted_onchip_memory2_3_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_0_instruction_master_readdatavalid = cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1 |
    cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1 |
    cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1 |
    cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_0_instruction_master_readdatavalid = cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    (cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in & dbs_counter_overflow) |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid;

  //cpu_0/instruction_master readdata mux, which is an e_mux
  assign cpu_0_instruction_master_readdata = ({32 {~(cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module & cpu_0_instruction_master_read)}} | cpu_0_jtag_debug_module_readdata_from_sa) &
    ({32 {~(cpu_0_instruction_master_qualified_request_nios_system_clock_2_in & cpu_0_instruction_master_read)}} | {nios_system_clock_2_in_readdata_from_sa[15 : 0],
    dbs_16_reg_segment_0}) &
    ({32 {~cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1}} | onchip_memory2_0_s1_readdata_from_sa) &
    ({32 {~cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1}} | onchip_memory2_1_s1_readdata_from_sa) &
    ({32 {~cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1}} | onchip_memory2_2_s1_readdata_from_sa) &
    ({32 {~cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1}} | onchip_memory2_3_s1_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_0_instruction_master_waitrequest = ~cpu_0_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_latency_counter <= 0;
      else 
        cpu_0_instruction_master_latency_counter <= p1_cpu_0_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_0_instruction_master_latency_counter = ((cpu_0_instruction_master_run & cpu_0_instruction_master_read))? latency_load_value :
    (cpu_0_instruction_master_latency_counter)? cpu_0_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({1 {cpu_0_instruction_master_requests_onchip_memory2_0_s1}} & 1) |
    ({1 {cpu_0_instruction_master_requests_onchip_memory2_1_s1}} & 1) |
    ({1 {cpu_0_instruction_master_requests_onchip_memory2_2_s1}} & 1) |
    ({1 {cpu_0_instruction_master_requests_onchip_memory2_3_s1}} & 1);

  //input to dbs-16 stored 0, which is an e_mux
  assign p1_dbs_16_reg_segment_0 = nios_system_clock_2_in_readdata_from_sa;

  //dbs register for dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_16_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_0_instruction_master_dbs_address[1]) == 0))
          dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
    end


  //dbs count increment, which is an e_mux
  assign cpu_0_instruction_master_dbs_increment = (cpu_0_instruction_master_requests_nios_system_clock_2_in)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_0_instruction_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_0_instruction_master_dbs_address + cpu_0_instruction_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_0_instruction_master_dbs_address <= next_dbs_address;
    end


  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = cpu_0_instruction_master_granted_nios_system_clock_2_in & cpu_0_instruction_master_read & 1 & 1 & ~nios_system_clock_2_in_waitrequest_from_sa;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_0_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_address_last_time <= 0;
      else 
        cpu_0_instruction_master_address_last_time <= cpu_0_instruction_master_address;
    end


  //cpu_0/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_0_instruction_master_waitrequest & (cpu_0_instruction_master_read);
    end


  //cpu_0_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_instruction_master_address != cpu_0_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_0_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_0_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_read_last_time <= 0;
      else 
        cpu_0_instruction_master_read_last_time <= cpu_0_instruction_master_read;
    end


  //cpu_0_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_instruction_master_read != cpu_0_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_0_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_0_altera_nios_custom_instr_floating_point_inst_s1_arbitrator (
                                                                          // inputs:
                                                                           clk,
                                                                           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done,
                                                                           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result,
                                                                           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select,
                                                                           cpu_0_custom_instruction_master_multi_clk_en,
                                                                           cpu_0_custom_instruction_master_multi_dataa,
                                                                           cpu_0_custom_instruction_master_multi_datab,
                                                                           cpu_0_custom_instruction_master_multi_n,
                                                                           cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1,
                                                                           reset_n,

                                                                          // outputs:
                                                                           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_clk_en,
                                                                           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_dataa,
                                                                           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_datab,
                                                                           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa,
                                                                           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_n,
                                                                           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_reset,
                                                                           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa,
                                                                           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_start
                                                                        )
;

  output           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  output  [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  output  [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_datab;
  output           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  output  [  1: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_n;
  output           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_reset;
  output  [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  output           cpu_0_altera_nios_custom_instr_floating_point_inst_s1_start;
  input            clk;
  input            cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done;
  input   [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result;
  input            cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select;
  input            cpu_0_custom_instruction_master_multi_clk_en;
  input   [ 31: 0] cpu_0_custom_instruction_master_multi_dataa;
  input   [ 31: 0] cpu_0_custom_instruction_master_multi_datab;
  input   [  7: 0] cpu_0_custom_instruction_master_multi_n;
  input            cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1;
  input            reset_n;

  wire             cpu_0_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  wire    [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  wire    [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_datab;
  wire             cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  wire    [  1: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_n;
  wire             cpu_0_altera_nios_custom_instr_floating_point_inst_s1_reset;
  wire    [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  wire             cpu_0_altera_nios_custom_instr_floating_point_inst_s1_start;
  assign cpu_0_altera_nios_custom_instr_floating_point_inst_s1_clk_en = cpu_0_custom_instruction_master_multi_clk_en;
  assign cpu_0_altera_nios_custom_instr_floating_point_inst_s1_dataa = cpu_0_custom_instruction_master_multi_dataa;
  assign cpu_0_altera_nios_custom_instr_floating_point_inst_s1_datab = cpu_0_custom_instruction_master_multi_datab;
  assign cpu_0_altera_nios_custom_instr_floating_point_inst_s1_n = cpu_0_custom_instruction_master_multi_n;
  assign cpu_0_altera_nios_custom_instr_floating_point_inst_s1_start = cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1;
  //assign cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa = cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa = cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result;

  //assign cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa = cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa = cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done;

  //cpu_0_altera_nios_custom_instr_floating_point_inst/s1 local reset_n, which is an e_assign
  assign cpu_0_altera_nios_custom_instr_floating_point_inst_s1_reset = ~reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_1_jtag_debug_module_arbitrator (
                                            // inputs:
                                             clk,
                                             cpu_1_data_master_address_to_slave,
                                             cpu_1_data_master_byteenable,
                                             cpu_1_data_master_debugaccess,
                                             cpu_1_data_master_latency_counter,
                                             cpu_1_data_master_read,
                                             cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                             cpu_1_data_master_write,
                                             cpu_1_data_master_writedata,
                                             cpu_1_instruction_master_address_to_slave,
                                             cpu_1_instruction_master_latency_counter,
                                             cpu_1_instruction_master_read,
                                             cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                             cpu_1_jtag_debug_module_readdata,
                                             cpu_1_jtag_debug_module_resetrequest,
                                             reset_n,

                                            // outputs:
                                             cpu_1_data_master_granted_cpu_1_jtag_debug_module,
                                             cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module,
                                             cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module,
                                             cpu_1_data_master_requests_cpu_1_jtag_debug_module,
                                             cpu_1_instruction_master_granted_cpu_1_jtag_debug_module,
                                             cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module,
                                             cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module,
                                             cpu_1_instruction_master_requests_cpu_1_jtag_debug_module,
                                             cpu_1_jtag_debug_module_address,
                                             cpu_1_jtag_debug_module_begintransfer,
                                             cpu_1_jtag_debug_module_byteenable,
                                             cpu_1_jtag_debug_module_chipselect,
                                             cpu_1_jtag_debug_module_debugaccess,
                                             cpu_1_jtag_debug_module_readdata_from_sa,
                                             cpu_1_jtag_debug_module_resetrequest_from_sa,
                                             cpu_1_jtag_debug_module_write,
                                             cpu_1_jtag_debug_module_writedata,
                                             d1_cpu_1_jtag_debug_module_end_xfer
                                          )
;

  output           cpu_1_data_master_granted_cpu_1_jtag_debug_module;
  output           cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module;
  output           cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module;
  output           cpu_1_data_master_requests_cpu_1_jtag_debug_module;
  output           cpu_1_instruction_master_granted_cpu_1_jtag_debug_module;
  output           cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module;
  output           cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module;
  output           cpu_1_instruction_master_requests_cpu_1_jtag_debug_module;
  output  [  8: 0] cpu_1_jtag_debug_module_address;
  output           cpu_1_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_1_jtag_debug_module_byteenable;
  output           cpu_1_jtag_debug_module_chipselect;
  output           cpu_1_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_1_jtag_debug_module_readdata_from_sa;
  output           cpu_1_jtag_debug_module_resetrequest_from_sa;
  output           cpu_1_jtag_debug_module_write;
  output  [ 31: 0] cpu_1_jtag_debug_module_writedata;
  output           d1_cpu_1_jtag_debug_module_end_xfer;
  input            clk;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input   [  3: 0] cpu_1_data_master_byteenable;
  input            cpu_1_data_master_debugaccess;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_1_instruction_master_address_to_slave;
  input            cpu_1_instruction_master_latency_counter;
  input            cpu_1_instruction_master_read;
  input            cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 31: 0] cpu_1_jtag_debug_module_readdata;
  input            cpu_1_jtag_debug_module_resetrequest;
  input            reset_n;

  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_cpu_1_jtag_debug_module;
  wire             cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module;
  wire             cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module;
  wire             cpu_1_data_master_requests_cpu_1_jtag_debug_module;
  wire             cpu_1_data_master_saved_grant_cpu_1_jtag_debug_module;
  wire             cpu_1_instruction_master_arbiterlock;
  wire             cpu_1_instruction_master_arbiterlock2;
  wire             cpu_1_instruction_master_continuerequest;
  wire             cpu_1_instruction_master_granted_cpu_1_jtag_debug_module;
  wire             cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module;
  wire             cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module;
  wire             cpu_1_instruction_master_requests_cpu_1_jtag_debug_module;
  wire             cpu_1_instruction_master_saved_grant_cpu_1_jtag_debug_module;
  wire    [  8: 0] cpu_1_jtag_debug_module_address;
  wire             cpu_1_jtag_debug_module_allgrants;
  wire             cpu_1_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_1_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_1_jtag_debug_module_any_continuerequest;
  reg     [  1: 0] cpu_1_jtag_debug_module_arb_addend;
  wire             cpu_1_jtag_debug_module_arb_counter_enable;
  reg     [  2: 0] cpu_1_jtag_debug_module_arb_share_counter;
  wire    [  2: 0] cpu_1_jtag_debug_module_arb_share_counter_next_value;
  wire    [  2: 0] cpu_1_jtag_debug_module_arb_share_set_values;
  wire    [  1: 0] cpu_1_jtag_debug_module_arb_winner;
  wire             cpu_1_jtag_debug_module_arbitration_holdoff_internal;
  wire             cpu_1_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_1_jtag_debug_module_begins_xfer;
  wire             cpu_1_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_1_jtag_debug_module_byteenable;
  wire             cpu_1_jtag_debug_module_chipselect;
  wire    [  3: 0] cpu_1_jtag_debug_module_chosen_master_double_vector;
  wire    [  1: 0] cpu_1_jtag_debug_module_chosen_master_rot_left;
  wire             cpu_1_jtag_debug_module_debugaccess;
  wire             cpu_1_jtag_debug_module_end_xfer;
  wire             cpu_1_jtag_debug_module_firsttransfer;
  wire    [  1: 0] cpu_1_jtag_debug_module_grant_vector;
  wire             cpu_1_jtag_debug_module_in_a_read_cycle;
  wire             cpu_1_jtag_debug_module_in_a_write_cycle;
  wire    [  1: 0] cpu_1_jtag_debug_module_master_qreq_vector;
  wire             cpu_1_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_1_jtag_debug_module_readdata_from_sa;
  reg              cpu_1_jtag_debug_module_reg_firsttransfer;
  wire             cpu_1_jtag_debug_module_resetrequest_from_sa;
  reg     [  1: 0] cpu_1_jtag_debug_module_saved_chosen_master_vector;
  reg              cpu_1_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_1_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_1_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_1_jtag_debug_module_waits_for_read;
  wire             cpu_1_jtag_debug_module_waits_for_write;
  wire             cpu_1_jtag_debug_module_write;
  wire    [ 31: 0] cpu_1_jtag_debug_module_writedata;
  reg              d1_cpu_1_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_1_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_1_data_master_granted_slave_cpu_1_jtag_debug_module;
  reg              last_cycle_cpu_1_instruction_master_granted_slave_cpu_1_jtag_debug_module;
  wire    [ 24: 0] shifted_address_to_cpu_1_jtag_debug_module_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_cpu_1_jtag_debug_module_from_cpu_1_instruction_master;
  wire             wait_for_cpu_1_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_1_jtag_debug_module_end_xfer;
    end


  assign cpu_1_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module | cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module));
  //assign cpu_1_jtag_debug_module_readdata_from_sa = cpu_1_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_1_jtag_debug_module_readdata_from_sa = cpu_1_jtag_debug_module_readdata;

  assign cpu_1_data_master_requests_cpu_1_jtag_debug_module = ({cpu_1_data_master_address_to_slave[24 : 11] , 11'b0} == 25'h1000) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //cpu_1_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_1_jtag_debug_module_arb_share_set_values = 1;

  //cpu_1_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_1_jtag_debug_module_non_bursting_master_requests = cpu_1_data_master_requests_cpu_1_jtag_debug_module |
    cpu_1_instruction_master_requests_cpu_1_jtag_debug_module |
    cpu_1_data_master_requests_cpu_1_jtag_debug_module |
    cpu_1_instruction_master_requests_cpu_1_jtag_debug_module;

  //cpu_1_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_1_jtag_debug_module_any_bursting_master_saved_grant = 0;

  //cpu_1_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_1_jtag_debug_module_arb_share_counter_next_value = cpu_1_jtag_debug_module_firsttransfer ? (cpu_1_jtag_debug_module_arb_share_set_values - 1) : |cpu_1_jtag_debug_module_arb_share_counter ? (cpu_1_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_1_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_1_jtag_debug_module_allgrants = (|cpu_1_jtag_debug_module_grant_vector) |
    (|cpu_1_jtag_debug_module_grant_vector) |
    (|cpu_1_jtag_debug_module_grant_vector) |
    (|cpu_1_jtag_debug_module_grant_vector);

  //cpu_1_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_1_jtag_debug_module_end_xfer = ~(cpu_1_jtag_debug_module_waits_for_read | cpu_1_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_1_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_1_jtag_debug_module = cpu_1_jtag_debug_module_end_xfer & (~cpu_1_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_1_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_1_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_1_jtag_debug_module & cpu_1_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_1_jtag_debug_module & ~cpu_1_jtag_debug_module_non_bursting_master_requests);

  //cpu_1_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_1_jtag_debug_module_arb_counter_enable)
          cpu_1_jtag_debug_module_arb_share_counter <= cpu_1_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_1_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_1_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_1_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_1_jtag_debug_module & ~cpu_1_jtag_debug_module_non_bursting_master_requests))
          cpu_1_jtag_debug_module_slavearbiterlockenable <= |cpu_1_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_1/data_master cpu_1/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = cpu_1_jtag_debug_module_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_1_jtag_debug_module_slavearbiterlockenable2 = |cpu_1_jtag_debug_module_arb_share_counter_next_value;

  //cpu_1/data_master cpu_1/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = cpu_1_jtag_debug_module_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/instruction_master cpu_1/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock = cpu_1_jtag_debug_module_slavearbiterlockenable & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master cpu_1/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock2 = cpu_1_jtag_debug_module_slavearbiterlockenable2 & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master granted cpu_1/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_instruction_master_granted_slave_cpu_1_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_1_instruction_master_granted_slave_cpu_1_jtag_debug_module <= cpu_1_instruction_master_saved_grant_cpu_1_jtag_debug_module ? 1 : (cpu_1_jtag_debug_module_arbitration_holdoff_internal | ~cpu_1_instruction_master_requests_cpu_1_jtag_debug_module) ? 0 : last_cycle_cpu_1_instruction_master_granted_slave_cpu_1_jtag_debug_module;
    end


  //cpu_1_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_1_instruction_master_continuerequest = last_cycle_cpu_1_instruction_master_granted_slave_cpu_1_jtag_debug_module & cpu_1_instruction_master_requests_cpu_1_jtag_debug_module;

  //cpu_1_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_1_jtag_debug_module_any_continuerequest = cpu_1_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest;

  assign cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module = cpu_1_data_master_requests_cpu_1_jtag_debug_module & ~((cpu_1_data_master_read & ((cpu_1_data_master_latency_counter != 0) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_1_instruction_master_arbiterlock);
  //local readdatavalid cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module, which is an e_mux
  assign cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module = cpu_1_data_master_granted_cpu_1_jtag_debug_module & cpu_1_data_master_read & ~cpu_1_jtag_debug_module_waits_for_read;

  //cpu_1_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_1_jtag_debug_module_writedata = cpu_1_data_master_writedata;

  assign cpu_1_instruction_master_requests_cpu_1_jtag_debug_module = (({cpu_1_instruction_master_address_to_slave[24 : 11] , 11'b0} == 25'h1000) & (cpu_1_instruction_master_read)) & cpu_1_instruction_master_read;
  //cpu_1/data_master granted cpu_1/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_cpu_1_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_cpu_1_jtag_debug_module <= cpu_1_data_master_saved_grant_cpu_1_jtag_debug_module ? 1 : (cpu_1_jtag_debug_module_arbitration_holdoff_internal | ~cpu_1_data_master_requests_cpu_1_jtag_debug_module) ? 0 : last_cycle_cpu_1_data_master_granted_slave_cpu_1_jtag_debug_module;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = last_cycle_cpu_1_data_master_granted_slave_cpu_1_jtag_debug_module & cpu_1_data_master_requests_cpu_1_jtag_debug_module;

  assign cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module = cpu_1_instruction_master_requests_cpu_1_jtag_debug_module & ~((cpu_1_instruction_master_read & ((cpu_1_instruction_master_latency_counter != 0) | (|cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_1_data_master_arbiterlock);
  //local readdatavalid cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module, which is an e_mux
  assign cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module = cpu_1_instruction_master_granted_cpu_1_jtag_debug_module & cpu_1_instruction_master_read & ~cpu_1_jtag_debug_module_waits_for_read;

  //allow new arb cycle for cpu_1/jtag_debug_module, which is an e_assign
  assign cpu_1_jtag_debug_module_allow_new_arb_cycle = ~cpu_1_data_master_arbiterlock & ~cpu_1_instruction_master_arbiterlock;

  //cpu_1/instruction_master assignment into master qualified-requests vector for cpu_1/jtag_debug_module, which is an e_assign
  assign cpu_1_jtag_debug_module_master_qreq_vector[0] = cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module;

  //cpu_1/instruction_master grant cpu_1/jtag_debug_module, which is an e_assign
  assign cpu_1_instruction_master_granted_cpu_1_jtag_debug_module = cpu_1_jtag_debug_module_grant_vector[0];

  //cpu_1/instruction_master saved-grant cpu_1/jtag_debug_module, which is an e_assign
  assign cpu_1_instruction_master_saved_grant_cpu_1_jtag_debug_module = cpu_1_jtag_debug_module_arb_winner[0] && cpu_1_instruction_master_requests_cpu_1_jtag_debug_module;

  //cpu_1/data_master assignment into master qualified-requests vector for cpu_1/jtag_debug_module, which is an e_assign
  assign cpu_1_jtag_debug_module_master_qreq_vector[1] = cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module;

  //cpu_1/data_master grant cpu_1/jtag_debug_module, which is an e_assign
  assign cpu_1_data_master_granted_cpu_1_jtag_debug_module = cpu_1_jtag_debug_module_grant_vector[1];

  //cpu_1/data_master saved-grant cpu_1/jtag_debug_module, which is an e_assign
  assign cpu_1_data_master_saved_grant_cpu_1_jtag_debug_module = cpu_1_jtag_debug_module_arb_winner[1] && cpu_1_data_master_requests_cpu_1_jtag_debug_module;

  //cpu_1/jtag_debug_module chosen-master double-vector, which is an e_assign
  assign cpu_1_jtag_debug_module_chosen_master_double_vector = {cpu_1_jtag_debug_module_master_qreq_vector, cpu_1_jtag_debug_module_master_qreq_vector} & ({~cpu_1_jtag_debug_module_master_qreq_vector, ~cpu_1_jtag_debug_module_master_qreq_vector} + cpu_1_jtag_debug_module_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_1_jtag_debug_module_arb_winner = (cpu_1_jtag_debug_module_allow_new_arb_cycle & | cpu_1_jtag_debug_module_grant_vector) ? cpu_1_jtag_debug_module_grant_vector : cpu_1_jtag_debug_module_saved_chosen_master_vector;

  //saved cpu_1_jtag_debug_module_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_jtag_debug_module_saved_chosen_master_vector <= 0;
      else if (cpu_1_jtag_debug_module_allow_new_arb_cycle)
          cpu_1_jtag_debug_module_saved_chosen_master_vector <= |cpu_1_jtag_debug_module_grant_vector ? cpu_1_jtag_debug_module_grant_vector : cpu_1_jtag_debug_module_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_1_jtag_debug_module_grant_vector = {(cpu_1_jtag_debug_module_chosen_master_double_vector[1] | cpu_1_jtag_debug_module_chosen_master_double_vector[3]),
    (cpu_1_jtag_debug_module_chosen_master_double_vector[0] | cpu_1_jtag_debug_module_chosen_master_double_vector[2])};

  //cpu_1/jtag_debug_module chosen master rotated left, which is an e_assign
  assign cpu_1_jtag_debug_module_chosen_master_rot_left = (cpu_1_jtag_debug_module_arb_winner << 1) ? (cpu_1_jtag_debug_module_arb_winner << 1) : 1;

  //cpu_1/jtag_debug_module's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_jtag_debug_module_arb_addend <= 1;
      else if (|cpu_1_jtag_debug_module_grant_vector)
          cpu_1_jtag_debug_module_arb_addend <= cpu_1_jtag_debug_module_end_xfer? cpu_1_jtag_debug_module_chosen_master_rot_left : cpu_1_jtag_debug_module_grant_vector;
    end


  assign cpu_1_jtag_debug_module_begintransfer = cpu_1_jtag_debug_module_begins_xfer;
  //assign cpu_1_jtag_debug_module_resetrequest_from_sa = cpu_1_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_1_jtag_debug_module_resetrequest_from_sa = cpu_1_jtag_debug_module_resetrequest;

  assign cpu_1_jtag_debug_module_chipselect = cpu_1_data_master_granted_cpu_1_jtag_debug_module | cpu_1_instruction_master_granted_cpu_1_jtag_debug_module;
  //cpu_1_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_1_jtag_debug_module_firsttransfer = cpu_1_jtag_debug_module_begins_xfer ? cpu_1_jtag_debug_module_unreg_firsttransfer : cpu_1_jtag_debug_module_reg_firsttransfer;

  //cpu_1_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_1_jtag_debug_module_unreg_firsttransfer = ~(cpu_1_jtag_debug_module_slavearbiterlockenable & cpu_1_jtag_debug_module_any_continuerequest);

  //cpu_1_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_1_jtag_debug_module_begins_xfer)
          cpu_1_jtag_debug_module_reg_firsttransfer <= cpu_1_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_1_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_1_jtag_debug_module_beginbursttransfer_internal = cpu_1_jtag_debug_module_begins_xfer;

  //cpu_1_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_1_jtag_debug_module_arbitration_holdoff_internal = cpu_1_jtag_debug_module_begins_xfer & cpu_1_jtag_debug_module_firsttransfer;

  //cpu_1_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_1_jtag_debug_module_write = cpu_1_data_master_granted_cpu_1_jtag_debug_module & cpu_1_data_master_write;

  assign shifted_address_to_cpu_1_jtag_debug_module_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  //cpu_1_jtag_debug_module_address mux, which is an e_mux
  assign cpu_1_jtag_debug_module_address = (cpu_1_data_master_granted_cpu_1_jtag_debug_module)? (shifted_address_to_cpu_1_jtag_debug_module_from_cpu_1_data_master >> 2) :
    (shifted_address_to_cpu_1_jtag_debug_module_from_cpu_1_instruction_master >> 2);

  assign shifted_address_to_cpu_1_jtag_debug_module_from_cpu_1_instruction_master = cpu_1_instruction_master_address_to_slave;
  //d1_cpu_1_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_1_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_1_jtag_debug_module_end_xfer <= cpu_1_jtag_debug_module_end_xfer;
    end


  //cpu_1_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_1_jtag_debug_module_waits_for_read = cpu_1_jtag_debug_module_in_a_read_cycle & cpu_1_jtag_debug_module_begins_xfer;

  //cpu_1_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_1_jtag_debug_module_in_a_read_cycle = (cpu_1_data_master_granted_cpu_1_jtag_debug_module & cpu_1_data_master_read) | (cpu_1_instruction_master_granted_cpu_1_jtag_debug_module & cpu_1_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_1_jtag_debug_module_in_a_read_cycle;

  //cpu_1_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_1_jtag_debug_module_waits_for_write = cpu_1_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_1_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_1_jtag_debug_module_in_a_write_cycle = cpu_1_data_master_granted_cpu_1_jtag_debug_module & cpu_1_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_1_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_1_jtag_debug_module_counter = 0;
  //cpu_1_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_1_jtag_debug_module_byteenable = (cpu_1_data_master_granted_cpu_1_jtag_debug_module)? cpu_1_data_master_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_1_jtag_debug_module_debugaccess = (cpu_1_data_master_granted_cpu_1_jtag_debug_module)? cpu_1_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_1/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_1_data_master_granted_cpu_1_jtag_debug_module + cpu_1_instruction_master_granted_cpu_1_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_1_data_master_saved_grant_cpu_1_jtag_debug_module + cpu_1_instruction_master_saved_grant_cpu_1_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_1_custom_instruction_master_arbitrator (
                                                    // inputs:
                                                     clk,
                                                     cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa,
                                                     cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa,
                                                     cpu_1_custom_instruction_master_multi_start,
                                                     reset_n,

                                                    // outputs:
                                                     cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select,
                                                     cpu_1_custom_instruction_master_multi_done,
                                                     cpu_1_custom_instruction_master_multi_result,
                                                     cpu_1_custom_instruction_master_reset_n,
                                                     cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1
                                                  )
;

  output           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select;
  output           cpu_1_custom_instruction_master_multi_done;
  output  [ 31: 0] cpu_1_custom_instruction_master_multi_result;
  output           cpu_1_custom_instruction_master_reset_n;
  output           cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1;
  input            clk;
  input            cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  input   [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  input            cpu_1_custom_instruction_master_multi_start;
  input            reset_n;

  wire             cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select;
  wire             cpu_1_custom_instruction_master_multi_done;
  wire    [ 31: 0] cpu_1_custom_instruction_master_multi_result;
  wire             cpu_1_custom_instruction_master_reset_n;
  wire             cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1;
  assign cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select = 1'b1;
  assign cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1 = cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select & cpu_1_custom_instruction_master_multi_start;
  //cpu_1_custom_instruction_master_multi_result mux, which is an e_mux
  assign cpu_1_custom_instruction_master_multi_result = {32 {cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select}} & cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;

  //multi_done mux, which is an e_mux
  assign cpu_1_custom_instruction_master_multi_done = {1 {cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select}} & cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;

  //cpu_1_custom_instruction_master_reset_n local reset_n, which is an e_assign
  assign cpu_1_custom_instruction_master_reset_n = reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_1_data_master_arbitrator (
                                      // inputs:
                                       clk,
                                       cpu_1_data_master_address,
                                       cpu_1_data_master_byteenable,
                                       cpu_1_data_master_byteenable_nios_system_clock_1_in,
                                       cpu_1_data_master_byteenable_nios_system_clock_8_in,
                                       cpu_1_data_master_byteenable_sram_0_avalon_sram_slave,
                                       cpu_1_data_master_granted_cpu_1_jtag_debug_module,
                                       cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave,
                                       cpu_1_data_master_granted_keys_s1,
                                       cpu_1_data_master_granted_mailbox_0_s1,
                                       cpu_1_data_master_granted_mailbox_1_s1,
                                       cpu_1_data_master_granted_mailbox_2_s1,
                                       cpu_1_data_master_granted_mailbox_3_s1,
                                       cpu_1_data_master_granted_nios_system_clock_1_in,
                                       cpu_1_data_master_granted_nios_system_clock_8_in,
                                       cpu_1_data_master_granted_onchip_memory2_0_s1,
                                       cpu_1_data_master_granted_onchip_memory2_1_s1,
                                       cpu_1_data_master_granted_onchip_memory2_2_s1,
                                       cpu_1_data_master_granted_onchip_memory2_3_s1,
                                       cpu_1_data_master_granted_performance_counter_0_control_slave,
                                       cpu_1_data_master_granted_sram_0_avalon_sram_slave,
                                       cpu_1_data_master_granted_sysid_control_slave,
                                       cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module,
                                       cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave,
                                       cpu_1_data_master_qualified_request_keys_s1,
                                       cpu_1_data_master_qualified_request_mailbox_0_s1,
                                       cpu_1_data_master_qualified_request_mailbox_1_s1,
                                       cpu_1_data_master_qualified_request_mailbox_2_s1,
                                       cpu_1_data_master_qualified_request_mailbox_3_s1,
                                       cpu_1_data_master_qualified_request_nios_system_clock_1_in,
                                       cpu_1_data_master_qualified_request_nios_system_clock_8_in,
                                       cpu_1_data_master_qualified_request_onchip_memory2_0_s1,
                                       cpu_1_data_master_qualified_request_onchip_memory2_1_s1,
                                       cpu_1_data_master_qualified_request_onchip_memory2_2_s1,
                                       cpu_1_data_master_qualified_request_onchip_memory2_3_s1,
                                       cpu_1_data_master_qualified_request_performance_counter_0_control_slave,
                                       cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave,
                                       cpu_1_data_master_qualified_request_sysid_control_slave,
                                       cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_1_data_master_read,
                                       cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module,
                                       cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave,
                                       cpu_1_data_master_read_data_valid_keys_s1,
                                       cpu_1_data_master_read_data_valid_mailbox_0_s1,
                                       cpu_1_data_master_read_data_valid_mailbox_1_s1,
                                       cpu_1_data_master_read_data_valid_mailbox_2_s1,
                                       cpu_1_data_master_read_data_valid_mailbox_3_s1,
                                       cpu_1_data_master_read_data_valid_nios_system_clock_1_in,
                                       cpu_1_data_master_read_data_valid_nios_system_clock_8_in,
                                       cpu_1_data_master_read_data_valid_onchip_memory2_0_s1,
                                       cpu_1_data_master_read_data_valid_onchip_memory2_1_s1,
                                       cpu_1_data_master_read_data_valid_onchip_memory2_2_s1,
                                       cpu_1_data_master_read_data_valid_onchip_memory2_3_s1,
                                       cpu_1_data_master_read_data_valid_performance_counter_0_control_slave,
                                       cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave,
                                       cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                       cpu_1_data_master_read_data_valid_sysid_control_slave,
                                       cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_1_data_master_requests_cpu_1_jtag_debug_module,
                                       cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave,
                                       cpu_1_data_master_requests_keys_s1,
                                       cpu_1_data_master_requests_mailbox_0_s1,
                                       cpu_1_data_master_requests_mailbox_1_s1,
                                       cpu_1_data_master_requests_mailbox_2_s1,
                                       cpu_1_data_master_requests_mailbox_3_s1,
                                       cpu_1_data_master_requests_nios_system_clock_1_in,
                                       cpu_1_data_master_requests_nios_system_clock_8_in,
                                       cpu_1_data_master_requests_onchip_memory2_0_s1,
                                       cpu_1_data_master_requests_onchip_memory2_1_s1,
                                       cpu_1_data_master_requests_onchip_memory2_2_s1,
                                       cpu_1_data_master_requests_onchip_memory2_3_s1,
                                       cpu_1_data_master_requests_performance_counter_0_control_slave,
                                       cpu_1_data_master_requests_sram_0_avalon_sram_slave,
                                       cpu_1_data_master_requests_sysid_control_slave,
                                       cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_1_data_master_write,
                                       cpu_1_data_master_writedata,
                                       cpu_1_jtag_debug_module_readdata_from_sa,
                                       d1_cpu_1_jtag_debug_module_end_xfer,
                                       d1_jtag_uart_1_avalon_jtag_slave_end_xfer,
                                       d1_keys_s1_end_xfer,
                                       d1_mailbox_0_s1_end_xfer,
                                       d1_mailbox_1_s1_end_xfer,
                                       d1_mailbox_2_s1_end_xfer,
                                       d1_mailbox_3_s1_end_xfer,
                                       d1_nios_system_clock_1_in_end_xfer,
                                       d1_nios_system_clock_8_in_end_xfer,
                                       d1_onchip_memory2_0_s1_end_xfer,
                                       d1_onchip_memory2_1_s1_end_xfer,
                                       d1_onchip_memory2_2_s1_end_xfer,
                                       d1_onchip_memory2_3_s1_end_xfer,
                                       d1_performance_counter_0_control_slave_end_xfer,
                                       d1_sram_0_avalon_sram_slave_end_xfer,
                                       d1_sysid_control_slave_end_xfer,
                                       d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer,
                                       jtag_uart_1_avalon_jtag_slave_irq_from_sa,
                                       jtag_uart_1_avalon_jtag_slave_readdata_from_sa,
                                       jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa,
                                       keys_s1_readdata_from_sa,
                                       mailbox_0_s1_readdata_from_sa,
                                       mailbox_1_s1_readdata_from_sa,
                                       mailbox_2_s1_readdata_from_sa,
                                       mailbox_3_s1_readdata_from_sa,
                                       nios_system_clock_1_in_readdata_from_sa,
                                       nios_system_clock_1_in_waitrequest_from_sa,
                                       nios_system_clock_8_in_readdata_from_sa,
                                       nios_system_clock_8_in_waitrequest_from_sa,
                                       onchip_memory2_0_s1_readdata_from_sa,
                                       onchip_memory2_1_s1_readdata_from_sa,
                                       onchip_memory2_2_s1_readdata_from_sa,
                                       onchip_memory2_3_s1_readdata_from_sa,
                                       performance_counter_0_control_slave_readdata_from_sa,
                                       reset_n,
                                       sram_0_avalon_sram_slave_readdata_from_sa,
                                       sysid_control_slave_readdata_from_sa,
                                       video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa,

                                      // outputs:
                                       cpu_1_data_master_address_to_slave,
                                       cpu_1_data_master_dbs_address,
                                       cpu_1_data_master_dbs_write_16,
                                       cpu_1_data_master_dbs_write_8,
                                       cpu_1_data_master_irq,
                                       cpu_1_data_master_latency_counter,
                                       cpu_1_data_master_readdata,
                                       cpu_1_data_master_readdatavalid,
                                       cpu_1_data_master_waitrequest
                                    )
;

  output  [ 24: 0] cpu_1_data_master_address_to_slave;
  output  [  1: 0] cpu_1_data_master_dbs_address;
  output  [ 15: 0] cpu_1_data_master_dbs_write_16;
  output  [  7: 0] cpu_1_data_master_dbs_write_8;
  output  [ 31: 0] cpu_1_data_master_irq;
  output           cpu_1_data_master_latency_counter;
  output  [ 31: 0] cpu_1_data_master_readdata;
  output           cpu_1_data_master_readdatavalid;
  output           cpu_1_data_master_waitrequest;
  input            clk;
  input   [ 24: 0] cpu_1_data_master_address;
  input   [  3: 0] cpu_1_data_master_byteenable;
  input   [  1: 0] cpu_1_data_master_byteenable_nios_system_clock_1_in;
  input            cpu_1_data_master_byteenable_nios_system_clock_8_in;
  input   [  1: 0] cpu_1_data_master_byteenable_sram_0_avalon_sram_slave;
  input            cpu_1_data_master_granted_cpu_1_jtag_debug_module;
  input            cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave;
  input            cpu_1_data_master_granted_keys_s1;
  input            cpu_1_data_master_granted_mailbox_0_s1;
  input            cpu_1_data_master_granted_mailbox_1_s1;
  input            cpu_1_data_master_granted_mailbox_2_s1;
  input            cpu_1_data_master_granted_mailbox_3_s1;
  input            cpu_1_data_master_granted_nios_system_clock_1_in;
  input            cpu_1_data_master_granted_nios_system_clock_8_in;
  input            cpu_1_data_master_granted_onchip_memory2_0_s1;
  input            cpu_1_data_master_granted_onchip_memory2_1_s1;
  input            cpu_1_data_master_granted_onchip_memory2_2_s1;
  input            cpu_1_data_master_granted_onchip_memory2_3_s1;
  input            cpu_1_data_master_granted_performance_counter_0_control_slave;
  input            cpu_1_data_master_granted_sram_0_avalon_sram_slave;
  input            cpu_1_data_master_granted_sysid_control_slave;
  input            cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module;
  input            cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave;
  input            cpu_1_data_master_qualified_request_keys_s1;
  input            cpu_1_data_master_qualified_request_mailbox_0_s1;
  input            cpu_1_data_master_qualified_request_mailbox_1_s1;
  input            cpu_1_data_master_qualified_request_mailbox_2_s1;
  input            cpu_1_data_master_qualified_request_mailbox_3_s1;
  input            cpu_1_data_master_qualified_request_nios_system_clock_1_in;
  input            cpu_1_data_master_qualified_request_nios_system_clock_8_in;
  input            cpu_1_data_master_qualified_request_onchip_memory2_0_s1;
  input            cpu_1_data_master_qualified_request_onchip_memory2_1_s1;
  input            cpu_1_data_master_qualified_request_onchip_memory2_2_s1;
  input            cpu_1_data_master_qualified_request_onchip_memory2_3_s1;
  input            cpu_1_data_master_qualified_request_performance_counter_0_control_slave;
  input            cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave;
  input            cpu_1_data_master_qualified_request_sysid_control_slave;
  input            cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module;
  input            cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave;
  input            cpu_1_data_master_read_data_valid_keys_s1;
  input            cpu_1_data_master_read_data_valid_mailbox_0_s1;
  input            cpu_1_data_master_read_data_valid_mailbox_1_s1;
  input            cpu_1_data_master_read_data_valid_mailbox_2_s1;
  input            cpu_1_data_master_read_data_valid_mailbox_3_s1;
  input            cpu_1_data_master_read_data_valid_nios_system_clock_1_in;
  input            cpu_1_data_master_read_data_valid_nios_system_clock_8_in;
  input            cpu_1_data_master_read_data_valid_onchip_memory2_0_s1;
  input            cpu_1_data_master_read_data_valid_onchip_memory2_1_s1;
  input            cpu_1_data_master_read_data_valid_onchip_memory2_2_s1;
  input            cpu_1_data_master_read_data_valid_onchip_memory2_3_s1;
  input            cpu_1_data_master_read_data_valid_performance_counter_0_control_slave;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_read_data_valid_sysid_control_slave;
  input            cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_1_data_master_requests_cpu_1_jtag_debug_module;
  input            cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave;
  input            cpu_1_data_master_requests_keys_s1;
  input            cpu_1_data_master_requests_mailbox_0_s1;
  input            cpu_1_data_master_requests_mailbox_1_s1;
  input            cpu_1_data_master_requests_mailbox_2_s1;
  input            cpu_1_data_master_requests_mailbox_3_s1;
  input            cpu_1_data_master_requests_nios_system_clock_1_in;
  input            cpu_1_data_master_requests_nios_system_clock_8_in;
  input            cpu_1_data_master_requests_onchip_memory2_0_s1;
  input            cpu_1_data_master_requests_onchip_memory2_1_s1;
  input            cpu_1_data_master_requests_onchip_memory2_2_s1;
  input            cpu_1_data_master_requests_onchip_memory2_3_s1;
  input            cpu_1_data_master_requests_performance_counter_0_control_slave;
  input            cpu_1_data_master_requests_sram_0_avalon_sram_slave;
  input            cpu_1_data_master_requests_sysid_control_slave;
  input            cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 31: 0] cpu_1_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_1_jtag_debug_module_end_xfer;
  input            d1_jtag_uart_1_avalon_jtag_slave_end_xfer;
  input            d1_keys_s1_end_xfer;
  input            d1_mailbox_0_s1_end_xfer;
  input            d1_mailbox_1_s1_end_xfer;
  input            d1_mailbox_2_s1_end_xfer;
  input            d1_mailbox_3_s1_end_xfer;
  input            d1_nios_system_clock_1_in_end_xfer;
  input            d1_nios_system_clock_8_in_end_xfer;
  input            d1_onchip_memory2_0_s1_end_xfer;
  input            d1_onchip_memory2_1_s1_end_xfer;
  input            d1_onchip_memory2_2_s1_end_xfer;
  input            d1_onchip_memory2_3_s1_end_xfer;
  input            d1_performance_counter_0_control_slave_end_xfer;
  input            d1_sram_0_avalon_sram_slave_end_xfer;
  input            d1_sysid_control_slave_end_xfer;
  input            d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer;
  input            jtag_uart_1_avalon_jtag_slave_irq_from_sa;
  input   [ 31: 0] jtag_uart_1_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa;
  input   [ 31: 0] keys_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_0_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_1_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_2_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_3_s1_readdata_from_sa;
  input   [ 15: 0] nios_system_clock_1_in_readdata_from_sa;
  input            nios_system_clock_1_in_waitrequest_from_sa;
  input   [  7: 0] nios_system_clock_8_in_readdata_from_sa;
  input            nios_system_clock_8_in_waitrequest_from_sa;
  input   [ 31: 0] onchip_memory2_0_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_1_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_2_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_3_s1_readdata_from_sa;
  input   [ 31: 0] performance_counter_0_control_slave_readdata_from_sa;
  input            reset_n;
  input   [ 15: 0] sram_0_avalon_sram_slave_readdata_from_sa;
  input   [ 31: 0] sysid_control_slave_readdata_from_sa;
  input   [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] cpu_1_data_master_address_last_time;
  wire    [ 24: 0] cpu_1_data_master_address_to_slave;
  reg     [  3: 0] cpu_1_data_master_byteenable_last_time;
  reg     [  1: 0] cpu_1_data_master_dbs_address;
  wire    [  1: 0] cpu_1_data_master_dbs_increment;
  reg     [  1: 0] cpu_1_data_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_1_data_master_dbs_rdv_counter_inc;
  wire    [ 15: 0] cpu_1_data_master_dbs_write_16;
  wire    [  7: 0] cpu_1_data_master_dbs_write_8;
  wire    [ 31: 0] cpu_1_data_master_irq;
  wire             cpu_1_data_master_is_granted_some_slave;
  reg              cpu_1_data_master_latency_counter;
  wire    [  1: 0] cpu_1_data_master_next_dbs_rdv_counter;
  reg              cpu_1_data_master_read_but_no_slave_selected;
  reg              cpu_1_data_master_read_last_time;
  wire    [ 31: 0] cpu_1_data_master_readdata;
  wire             cpu_1_data_master_readdatavalid;
  wire             cpu_1_data_master_run;
  wire             cpu_1_data_master_waitrequest;
  reg              cpu_1_data_master_write_last_time;
  reg     [ 31: 0] cpu_1_data_master_writedata_last_time;
  reg     [ 15: 0] dbs_16_reg_segment_0;
  reg     [  7: 0] dbs_8_reg_segment_0;
  reg     [  7: 0] dbs_8_reg_segment_1;
  reg     [  7: 0] dbs_8_reg_segment_2;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire             p1_cpu_1_data_master_latency_counter;
  wire    [ 15: 0] p1_dbs_16_reg_segment_0;
  wire    [  7: 0] p1_dbs_8_reg_segment_0;
  wire    [  7: 0] p1_dbs_8_reg_segment_1;
  wire    [  7: 0] p1_dbs_8_reg_segment_2;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_1_data_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  wire             r_3;
  wire             r_4;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module | ~cpu_1_data_master_requests_cpu_1_jtag_debug_module) & (cpu_1_data_master_granted_cpu_1_jtag_debug_module | ~cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module) & ((~cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module | ~cpu_1_data_master_read | (1 & ~d1_cpu_1_jtag_debug_module_end_xfer & cpu_1_data_master_read))) & ((~cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module | ~cpu_1_data_master_write | (1 & cpu_1_data_master_write))) & 1 & (cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave | ~cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave) & ((~cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & ~jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa & (cpu_1_data_master_read | cpu_1_data_master_write)))) & ((~cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & ~jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa & (cpu_1_data_master_read | cpu_1_data_master_write)))) & 1 & (cpu_1_data_master_qualified_request_keys_s1 | ~cpu_1_data_master_requests_keys_s1) & (cpu_1_data_master_granted_keys_s1 | ~cpu_1_data_master_qualified_request_keys_s1) & ((~cpu_1_data_master_qualified_request_keys_s1 | ~cpu_1_data_master_read | (1 & ~d1_keys_s1_end_xfer & cpu_1_data_master_read))) & ((~cpu_1_data_master_qualified_request_keys_s1 | ~cpu_1_data_master_write | (1 & cpu_1_data_master_write))) & 1 & (cpu_1_data_master_qualified_request_mailbox_0_s1 | ~cpu_1_data_master_requests_mailbox_0_s1) & (cpu_1_data_master_granted_mailbox_0_s1 | ~cpu_1_data_master_qualified_request_mailbox_0_s1) & ((~cpu_1_data_master_qualified_request_mailbox_0_s1 | ~cpu_1_data_master_read | (1 & ~d1_mailbox_0_s1_end_xfer & cpu_1_data_master_read))) & ((~cpu_1_data_master_qualified_request_mailbox_0_s1 | ~cpu_1_data_master_write | (1 & cpu_1_data_master_write)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_1_data_master_run = r_0 & r_1 & r_2 & r_3 & r_4;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_1_data_master_qualified_request_mailbox_1_s1 | ~cpu_1_data_master_requests_mailbox_1_s1) & (cpu_1_data_master_granted_mailbox_1_s1 | ~cpu_1_data_master_qualified_request_mailbox_1_s1) & ((~cpu_1_data_master_qualified_request_mailbox_1_s1 | ~cpu_1_data_master_read | (1 & ~d1_mailbox_1_s1_end_xfer & cpu_1_data_master_read))) & ((~cpu_1_data_master_qualified_request_mailbox_1_s1 | ~cpu_1_data_master_write | (1 & cpu_1_data_master_write))) & 1 & (cpu_1_data_master_qualified_request_mailbox_2_s1 | ~cpu_1_data_master_requests_mailbox_2_s1) & (cpu_1_data_master_granted_mailbox_2_s1 | ~cpu_1_data_master_qualified_request_mailbox_2_s1) & ((~cpu_1_data_master_qualified_request_mailbox_2_s1 | ~cpu_1_data_master_read | (1 & ~d1_mailbox_2_s1_end_xfer & cpu_1_data_master_read))) & ((~cpu_1_data_master_qualified_request_mailbox_2_s1 | ~cpu_1_data_master_write | (1 & cpu_1_data_master_write))) & 1 & (cpu_1_data_master_qualified_request_mailbox_3_s1 | ~cpu_1_data_master_requests_mailbox_3_s1) & (cpu_1_data_master_granted_mailbox_3_s1 | ~cpu_1_data_master_qualified_request_mailbox_3_s1) & ((~cpu_1_data_master_qualified_request_mailbox_3_s1 | ~cpu_1_data_master_read | (1 & ~d1_mailbox_3_s1_end_xfer & cpu_1_data_master_read))) & ((~cpu_1_data_master_qualified_request_mailbox_3_s1 | ~cpu_1_data_master_write | (1 & cpu_1_data_master_write))) & 1 & (cpu_1_data_master_qualified_request_nios_system_clock_1_in | (cpu_1_data_master_write & !cpu_1_data_master_byteenable_nios_system_clock_1_in & cpu_1_data_master_dbs_address[1]) | ~cpu_1_data_master_requests_nios_system_clock_1_in) & ((~cpu_1_data_master_qualified_request_nios_system_clock_1_in | ~cpu_1_data_master_read | (1 & ~nios_system_clock_1_in_waitrequest_from_sa & (cpu_1_data_master_dbs_address[1]) & cpu_1_data_master_read))) & ((~cpu_1_data_master_qualified_request_nios_system_clock_1_in | ~cpu_1_data_master_write | (1 & ~nios_system_clock_1_in_waitrequest_from_sa & (cpu_1_data_master_dbs_address[1]) & cpu_1_data_master_write)));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & ((cpu_1_data_master_qualified_request_nios_system_clock_8_in | ((cpu_1_data_master_write & !cpu_1_data_master_byteenable_nios_system_clock_8_in & cpu_1_data_master_dbs_address[1] & cpu_1_data_master_dbs_address[0])) | ~cpu_1_data_master_requests_nios_system_clock_8_in)) & ((~cpu_1_data_master_qualified_request_nios_system_clock_8_in | ~cpu_1_data_master_read | (1 & ~nios_system_clock_8_in_waitrequest_from_sa & (cpu_1_data_master_dbs_address[1] & cpu_1_data_master_dbs_address[0]) & cpu_1_data_master_read))) & ((~cpu_1_data_master_qualified_request_nios_system_clock_8_in | ~cpu_1_data_master_write | (1 & ~nios_system_clock_8_in_waitrequest_from_sa & (cpu_1_data_master_dbs_address[1] & cpu_1_data_master_dbs_address[0]) & cpu_1_data_master_write))) & 1 & (cpu_1_data_master_qualified_request_onchip_memory2_0_s1 | ~cpu_1_data_master_requests_onchip_memory2_0_s1) & (cpu_1_data_master_granted_onchip_memory2_0_s1 | ~cpu_1_data_master_qualified_request_onchip_memory2_0_s1) & ((~cpu_1_data_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write)))) & ((~cpu_1_data_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write)))) & 1 & (cpu_1_data_master_qualified_request_onchip_memory2_1_s1 | ~cpu_1_data_master_requests_onchip_memory2_1_s1) & (cpu_1_data_master_granted_onchip_memory2_1_s1 | ~cpu_1_data_master_qualified_request_onchip_memory2_1_s1) & ((~cpu_1_data_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write)))) & ((~cpu_1_data_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write)))) & 1 & (cpu_1_data_master_qualified_request_onchip_memory2_2_s1 | ~cpu_1_data_master_requests_onchip_memory2_2_s1) & (cpu_1_data_master_granted_onchip_memory2_2_s1 | ~cpu_1_data_master_qualified_request_onchip_memory2_2_s1) & ((~cpu_1_data_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write)))) & ((~cpu_1_data_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write))));

  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (cpu_1_data_master_qualified_request_onchip_memory2_3_s1 | ~cpu_1_data_master_requests_onchip_memory2_3_s1) & (cpu_1_data_master_granted_onchip_memory2_3_s1 | ~cpu_1_data_master_qualified_request_onchip_memory2_3_s1) & ((~cpu_1_data_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write)))) & ((~cpu_1_data_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write)))) & 1 & (cpu_1_data_master_qualified_request_performance_counter_0_control_slave | ~cpu_1_data_master_requests_performance_counter_0_control_slave) & (cpu_1_data_master_granted_performance_counter_0_control_slave | ~cpu_1_data_master_qualified_request_performance_counter_0_control_slave) & ((~cpu_1_data_master_qualified_request_performance_counter_0_control_slave | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write)))) & ((~cpu_1_data_master_qualified_request_performance_counter_0_control_slave | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write)))) & 1 & (cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave | (cpu_1_data_master_write & !cpu_1_data_master_byteenable_sram_0_avalon_sram_slave & cpu_1_data_master_dbs_address[1]) | ~cpu_1_data_master_requests_sram_0_avalon_sram_slave) & (cpu_1_data_master_granted_sram_0_avalon_sram_slave | ~cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave) & ((~cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_1_data_master_read | (1 & (cpu_1_data_master_dbs_address[1]) & cpu_1_data_master_read))) & ((~cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_1_data_master_write | (1 & (cpu_1_data_master_dbs_address[1]) & cpu_1_data_master_write))) & 1 & (cpu_1_data_master_qualified_request_sysid_control_slave | ~cpu_1_data_master_requests_sysid_control_slave) & (cpu_1_data_master_granted_sysid_control_slave | ~cpu_1_data_master_qualified_request_sysid_control_slave) & ((~cpu_1_data_master_qualified_request_sysid_control_slave | ~cpu_1_data_master_read | (1 & ~d1_sysid_control_slave_end_xfer & cpu_1_data_master_read))) & ((~cpu_1_data_master_qualified_request_sysid_control_slave | ~cpu_1_data_master_write | (1 & cpu_1_data_master_write)));

  //r_4 master_run cascaded wait assignment, which is an e_assign
  assign r_4 = 1 & (cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) & (cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave | ~cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave) & ((~cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write)))) & ((~cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~(cpu_1_data_master_read | cpu_1_data_master_write) | (1 & (cpu_1_data_master_read | cpu_1_data_master_write))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_1_data_master_address_to_slave = cpu_1_data_master_address[24 : 0];

  //cpu_1_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_read_but_no_slave_selected <= 0;
      else 
        cpu_1_data_master_read_but_no_slave_selected <= cpu_1_data_master_read & cpu_1_data_master_run & ~cpu_1_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_1_data_master_is_granted_some_slave = cpu_1_data_master_granted_cpu_1_jtag_debug_module |
    cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave |
    cpu_1_data_master_granted_keys_s1 |
    cpu_1_data_master_granted_mailbox_0_s1 |
    cpu_1_data_master_granted_mailbox_1_s1 |
    cpu_1_data_master_granted_mailbox_2_s1 |
    cpu_1_data_master_granted_mailbox_3_s1 |
    cpu_1_data_master_granted_nios_system_clock_1_in |
    cpu_1_data_master_granted_nios_system_clock_8_in |
    cpu_1_data_master_granted_onchip_memory2_0_s1 |
    cpu_1_data_master_granted_onchip_memory2_1_s1 |
    cpu_1_data_master_granted_onchip_memory2_2_s1 |
    cpu_1_data_master_granted_onchip_memory2_3_s1 |
    cpu_1_data_master_granted_performance_counter_0_control_slave |
    cpu_1_data_master_granted_sram_0_avalon_sram_slave |
    cpu_1_data_master_granted_sysid_control_slave |
    cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_1_data_master_readdatavalid = cpu_1_data_master_read_data_valid_onchip_memory2_0_s1 |
    cpu_1_data_master_read_data_valid_onchip_memory2_1_s1 |
    cpu_1_data_master_read_data_valid_onchip_memory2_2_s1 |
    cpu_1_data_master_read_data_valid_onchip_memory2_3_s1 |
    cpu_1_data_master_read_data_valid_performance_counter_0_control_slave |
    (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave & dbs_rdv_counter_overflow) |
    cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_1_data_master_readdatavalid = cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_data_valid_keys_s1 |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_data_valid_mailbox_0_s1 |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_data_valid_mailbox_1_s1 |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_data_valid_mailbox_2_s1 |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_data_valid_mailbox_3_s1 |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    (cpu_1_data_master_read_data_valid_nios_system_clock_1_in & dbs_counter_overflow) |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    (cpu_1_data_master_read_data_valid_nios_system_clock_8_in & dbs_counter_overflow) |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid |
    cpu_1_data_master_read_data_valid_sysid_control_slave |
    cpu_1_data_master_read_but_no_slave_selected |
    pre_flush_cpu_1_data_master_readdatavalid;

  //cpu_1/data_master readdata mux, which is an e_mux
  assign cpu_1_data_master_readdata = ({32 {~(cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module & cpu_1_data_master_read)}} | cpu_1_jtag_debug_module_readdata_from_sa) &
    ({32 {~(cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave & cpu_1_data_master_read)}} | jtag_uart_1_avalon_jtag_slave_readdata_from_sa) &
    ({32 {~(cpu_1_data_master_qualified_request_keys_s1 & cpu_1_data_master_read)}} | keys_s1_readdata_from_sa) &
    ({32 {~(cpu_1_data_master_qualified_request_mailbox_0_s1 & cpu_1_data_master_read)}} | mailbox_0_s1_readdata_from_sa) &
    ({32 {~(cpu_1_data_master_qualified_request_mailbox_1_s1 & cpu_1_data_master_read)}} | mailbox_1_s1_readdata_from_sa) &
    ({32 {~(cpu_1_data_master_qualified_request_mailbox_2_s1 & cpu_1_data_master_read)}} | mailbox_2_s1_readdata_from_sa) &
    ({32 {~(cpu_1_data_master_qualified_request_mailbox_3_s1 & cpu_1_data_master_read)}} | mailbox_3_s1_readdata_from_sa) &
    ({32 {~(cpu_1_data_master_qualified_request_nios_system_clock_1_in & cpu_1_data_master_read)}} | {nios_system_clock_1_in_readdata_from_sa[15 : 0],
    dbs_16_reg_segment_0}) &
    ({32 {~(cpu_1_data_master_qualified_request_nios_system_clock_8_in & cpu_1_data_master_read)}} | {nios_system_clock_8_in_readdata_from_sa[7 : 0],
    dbs_8_reg_segment_2,
    dbs_8_reg_segment_1,
    dbs_8_reg_segment_0}) &
    ({32 {~cpu_1_data_master_read_data_valid_onchip_memory2_0_s1}} | onchip_memory2_0_s1_readdata_from_sa) &
    ({32 {~cpu_1_data_master_read_data_valid_onchip_memory2_1_s1}} | onchip_memory2_1_s1_readdata_from_sa) &
    ({32 {~cpu_1_data_master_read_data_valid_onchip_memory2_2_s1}} | onchip_memory2_2_s1_readdata_from_sa) &
    ({32 {~cpu_1_data_master_read_data_valid_onchip_memory2_3_s1}} | onchip_memory2_3_s1_readdata_from_sa) &
    ({32 {~cpu_1_data_master_read_data_valid_performance_counter_0_control_slave}} | performance_counter_0_control_slave_readdata_from_sa) &
    ({32 {~cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave}} | {sram_0_avalon_sram_slave_readdata_from_sa[15 : 0],
    dbs_latent_16_reg_segment_0}) &
    ({32 {~(cpu_1_data_master_qualified_request_sysid_control_slave & cpu_1_data_master_read)}} | sysid_control_slave_readdata_from_sa) &
    ({32 {~cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave}} | video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_1_data_master_waitrequest = ~cpu_1_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_latency_counter <= 0;
      else 
        cpu_1_data_master_latency_counter <= p1_cpu_1_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_1_data_master_latency_counter = ((cpu_1_data_master_run & cpu_1_data_master_read))? latency_load_value :
    (cpu_1_data_master_latency_counter)? cpu_1_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({1 {cpu_1_data_master_requests_onchip_memory2_0_s1}} & 1) |
    ({1 {cpu_1_data_master_requests_onchip_memory2_1_s1}} & 1) |
    ({1 {cpu_1_data_master_requests_onchip_memory2_2_s1}} & 1) |
    ({1 {cpu_1_data_master_requests_onchip_memory2_3_s1}} & 1) |
    ({1 {cpu_1_data_master_requests_performance_counter_0_control_slave}} & 1) |
    ({1 {cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave}} & 1);

  //irq assign, which is an e_assign
  assign cpu_1_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    jtag_uart_1_avalon_jtag_slave_irq_from_sa,
    1'b0};

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (((~0) & cpu_1_data_master_requests_nios_system_clock_1_in & cpu_1_data_master_write & !cpu_1_data_master_byteenable_nios_system_clock_1_in)) |
    (cpu_1_data_master_granted_nios_system_clock_1_in & cpu_1_data_master_read & 1 & 1 & ~nios_system_clock_1_in_waitrequest_from_sa) |
    (cpu_1_data_master_granted_nios_system_clock_1_in & cpu_1_data_master_write & 1 & 1 & ~nios_system_clock_1_in_waitrequest_from_sa) |
    (((~0) & cpu_1_data_master_requests_nios_system_clock_8_in & cpu_1_data_master_write & !cpu_1_data_master_byteenable_nios_system_clock_8_in)) |
    (cpu_1_data_master_granted_nios_system_clock_8_in & cpu_1_data_master_read & 1 & 1 & ~nios_system_clock_8_in_waitrequest_from_sa) |
    (cpu_1_data_master_granted_nios_system_clock_8_in & cpu_1_data_master_write & 1 & 1 & ~nios_system_clock_8_in_waitrequest_from_sa) |
    (((~0) & cpu_1_data_master_requests_sram_0_avalon_sram_slave & cpu_1_data_master_write & !cpu_1_data_master_byteenable_sram_0_avalon_sram_slave)) |
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave & cpu_1_data_master_read & 1 & 1) |
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave & cpu_1_data_master_write & 1 & 1);

  //input to dbs-16 stored 0, which is an e_mux
  assign p1_dbs_16_reg_segment_0 = nios_system_clock_1_in_readdata_from_sa;

  //dbs register for dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_16_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_1_data_master_dbs_address[1]) == 0))
          dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
    end


  //mux write dbs 1, which is an e_mux
  assign cpu_1_data_master_dbs_write_16 = (cpu_1_data_master_dbs_address[1])? cpu_1_data_master_writedata[31 : 16] :
    (~(cpu_1_data_master_dbs_address[1]))? cpu_1_data_master_writedata[15 : 0] :
    (cpu_1_data_master_dbs_address[1])? cpu_1_data_master_writedata[31 : 16] :
    cpu_1_data_master_writedata[15 : 0];

  //dbs count increment, which is an e_mux
  assign cpu_1_data_master_dbs_increment = (cpu_1_data_master_requests_nios_system_clock_1_in)? 2 :
    (cpu_1_data_master_requests_nios_system_clock_8_in)? 1 :
    (cpu_1_data_master_requests_sram_0_avalon_sram_slave)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_1_data_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_1_data_master_dbs_address + cpu_1_data_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_1_data_master_dbs_address <= next_dbs_address;
    end


  //input to dbs-8 stored 0, which is an e_mux
  assign p1_dbs_8_reg_segment_0 = nios_system_clock_8_in_readdata_from_sa;

  //dbs register for dbs-8 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_1_data_master_dbs_address[1 : 0]) == 0))
          dbs_8_reg_segment_0 <= p1_dbs_8_reg_segment_0;
    end


  //input to dbs-8 stored 1, which is an e_mux
  assign p1_dbs_8_reg_segment_1 = nios_system_clock_8_in_readdata_from_sa;

  //dbs register for dbs-8 segment 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_1 <= 0;
      else if (dbs_count_enable & ((cpu_1_data_master_dbs_address[1 : 0]) == 1))
          dbs_8_reg_segment_1 <= p1_dbs_8_reg_segment_1;
    end


  //input to dbs-8 stored 2, which is an e_mux
  assign p1_dbs_8_reg_segment_2 = nios_system_clock_8_in_readdata_from_sa;

  //dbs register for dbs-8 segment 2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_2 <= 0;
      else if (dbs_count_enable & ((cpu_1_data_master_dbs_address[1 : 0]) == 2))
          dbs_8_reg_segment_2 <= p1_dbs_8_reg_segment_2;
    end


  //mux write dbs 2, which is an e_mux
  assign cpu_1_data_master_dbs_write_8 = ((cpu_1_data_master_dbs_address[1 : 0] == 0))? cpu_1_data_master_writedata[7 : 0] :
    ((cpu_1_data_master_dbs_address[1 : 0] == 1))? cpu_1_data_master_writedata[15 : 8] :
    ((cpu_1_data_master_dbs_address[1 : 0] == 2))? cpu_1_data_master_writedata[23 : 16] :
    cpu_1_data_master_writedata[31 : 24];

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = sram_0_avalon_sram_slave_readdata_from_sa;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_1_data_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_1_data_master_next_dbs_rdv_counter = cpu_1_data_master_dbs_rdv_counter + cpu_1_data_master_dbs_rdv_counter_inc;

  //cpu_1_data_master_rdv_inc_mux, which is an e_mux
  assign cpu_1_data_master_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_1_data_master_dbs_rdv_counter <= cpu_1_data_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_1_data_master_dbs_rdv_counter[1] & ~cpu_1_data_master_next_dbs_rdv_counter[1];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_1_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_address_last_time <= 0;
      else 
        cpu_1_data_master_address_last_time <= cpu_1_data_master_address;
    end


  //cpu_1/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_1_data_master_waitrequest & (cpu_1_data_master_read | cpu_1_data_master_write);
    end


  //cpu_1_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_1_data_master_address != cpu_1_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_1_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_1_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_byteenable_last_time <= 0;
      else 
        cpu_1_data_master_byteenable_last_time <= cpu_1_data_master_byteenable;
    end


  //cpu_1_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_1_data_master_byteenable != cpu_1_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_1_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_1_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_read_last_time <= 0;
      else 
        cpu_1_data_master_read_last_time <= cpu_1_data_master_read;
    end


  //cpu_1_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_1_data_master_read != cpu_1_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_1_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_1_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_write_last_time <= 0;
      else 
        cpu_1_data_master_write_last_time <= cpu_1_data_master_write;
    end


  //cpu_1_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_1_data_master_write != cpu_1_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_1_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_1_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_writedata_last_time <= 0;
      else 
        cpu_1_data_master_writedata_last_time <= cpu_1_data_master_writedata;
    end


  //cpu_1_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_1_data_master_writedata != cpu_1_data_master_writedata_last_time) & cpu_1_data_master_write)
        begin
          $write("%0d ns: cpu_1_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_1_instruction_master_arbitrator (
                                             // inputs:
                                              clk,
                                              cpu_1_instruction_master_address,
                                              cpu_1_instruction_master_granted_cpu_1_jtag_debug_module,
                                              cpu_1_instruction_master_granted_nios_system_clock_0_in,
                                              cpu_1_instruction_master_granted_onchip_memory2_0_s1,
                                              cpu_1_instruction_master_granted_onchip_memory2_1_s1,
                                              cpu_1_instruction_master_granted_onchip_memory2_2_s1,
                                              cpu_1_instruction_master_granted_onchip_memory2_3_s1,
                                              cpu_1_instruction_master_granted_sram_0_avalon_sram_slave,
                                              cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module,
                                              cpu_1_instruction_master_qualified_request_nios_system_clock_0_in,
                                              cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1,
                                              cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1,
                                              cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1,
                                              cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1,
                                              cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave,
                                              cpu_1_instruction_master_read,
                                              cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module,
                                              cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in,
                                              cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1,
                                              cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1,
                                              cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1,
                                              cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1,
                                              cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave,
                                              cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                              cpu_1_instruction_master_requests_cpu_1_jtag_debug_module,
                                              cpu_1_instruction_master_requests_nios_system_clock_0_in,
                                              cpu_1_instruction_master_requests_onchip_memory2_0_s1,
                                              cpu_1_instruction_master_requests_onchip_memory2_1_s1,
                                              cpu_1_instruction_master_requests_onchip_memory2_2_s1,
                                              cpu_1_instruction_master_requests_onchip_memory2_3_s1,
                                              cpu_1_instruction_master_requests_sram_0_avalon_sram_slave,
                                              cpu_1_jtag_debug_module_readdata_from_sa,
                                              d1_cpu_1_jtag_debug_module_end_xfer,
                                              d1_nios_system_clock_0_in_end_xfer,
                                              d1_onchip_memory2_0_s1_end_xfer,
                                              d1_onchip_memory2_1_s1_end_xfer,
                                              d1_onchip_memory2_2_s1_end_xfer,
                                              d1_onchip_memory2_3_s1_end_xfer,
                                              d1_sram_0_avalon_sram_slave_end_xfer,
                                              nios_system_clock_0_in_readdata_from_sa,
                                              nios_system_clock_0_in_waitrequest_from_sa,
                                              onchip_memory2_0_s1_readdata_from_sa,
                                              onchip_memory2_1_s1_readdata_from_sa,
                                              onchip_memory2_2_s1_readdata_from_sa,
                                              onchip_memory2_3_s1_readdata_from_sa,
                                              reset_n,
                                              sram_0_avalon_sram_slave_readdata_from_sa,

                                             // outputs:
                                              cpu_1_instruction_master_address_to_slave,
                                              cpu_1_instruction_master_dbs_address,
                                              cpu_1_instruction_master_latency_counter,
                                              cpu_1_instruction_master_readdata,
                                              cpu_1_instruction_master_readdatavalid,
                                              cpu_1_instruction_master_waitrequest
                                           )
;

  output  [ 24: 0] cpu_1_instruction_master_address_to_slave;
  output  [  1: 0] cpu_1_instruction_master_dbs_address;
  output           cpu_1_instruction_master_latency_counter;
  output  [ 31: 0] cpu_1_instruction_master_readdata;
  output           cpu_1_instruction_master_readdatavalid;
  output           cpu_1_instruction_master_waitrequest;
  input            clk;
  input   [ 24: 0] cpu_1_instruction_master_address;
  input            cpu_1_instruction_master_granted_cpu_1_jtag_debug_module;
  input            cpu_1_instruction_master_granted_nios_system_clock_0_in;
  input            cpu_1_instruction_master_granted_onchip_memory2_0_s1;
  input            cpu_1_instruction_master_granted_onchip_memory2_1_s1;
  input            cpu_1_instruction_master_granted_onchip_memory2_2_s1;
  input            cpu_1_instruction_master_granted_onchip_memory2_3_s1;
  input            cpu_1_instruction_master_granted_sram_0_avalon_sram_slave;
  input            cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module;
  input            cpu_1_instruction_master_qualified_request_nios_system_clock_0_in;
  input            cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1;
  input            cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1;
  input            cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1;
  input            cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1;
  input            cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  input            cpu_1_instruction_master_read;
  input            cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module;
  input            cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in;
  input            cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1;
  input            cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1;
  input            cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1;
  input            cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1;
  input            cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  input            cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_instruction_master_requests_cpu_1_jtag_debug_module;
  input            cpu_1_instruction_master_requests_nios_system_clock_0_in;
  input            cpu_1_instruction_master_requests_onchip_memory2_0_s1;
  input            cpu_1_instruction_master_requests_onchip_memory2_1_s1;
  input            cpu_1_instruction_master_requests_onchip_memory2_2_s1;
  input            cpu_1_instruction_master_requests_onchip_memory2_3_s1;
  input            cpu_1_instruction_master_requests_sram_0_avalon_sram_slave;
  input   [ 31: 0] cpu_1_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_1_jtag_debug_module_end_xfer;
  input            d1_nios_system_clock_0_in_end_xfer;
  input            d1_onchip_memory2_0_s1_end_xfer;
  input            d1_onchip_memory2_1_s1_end_xfer;
  input            d1_onchip_memory2_2_s1_end_xfer;
  input            d1_onchip_memory2_3_s1_end_xfer;
  input            d1_sram_0_avalon_sram_slave_end_xfer;
  input   [ 15: 0] nios_system_clock_0_in_readdata_from_sa;
  input            nios_system_clock_0_in_waitrequest_from_sa;
  input   [ 31: 0] onchip_memory2_0_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_1_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_2_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_3_s1_readdata_from_sa;
  input            reset_n;
  input   [ 15: 0] sram_0_avalon_sram_slave_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] cpu_1_instruction_master_address_last_time;
  wire    [ 24: 0] cpu_1_instruction_master_address_to_slave;
  reg     [  1: 0] cpu_1_instruction_master_dbs_address;
  wire    [  1: 0] cpu_1_instruction_master_dbs_increment;
  reg     [  1: 0] cpu_1_instruction_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_1_instruction_master_dbs_rdv_counter_inc;
  wire             cpu_1_instruction_master_is_granted_some_slave;
  reg              cpu_1_instruction_master_latency_counter;
  wire    [  1: 0] cpu_1_instruction_master_next_dbs_rdv_counter;
  reg              cpu_1_instruction_master_read_but_no_slave_selected;
  reg              cpu_1_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_1_instruction_master_readdata;
  wire             cpu_1_instruction_master_readdatavalid;
  wire             cpu_1_instruction_master_run;
  wire             cpu_1_instruction_master_waitrequest;
  reg     [ 15: 0] dbs_16_reg_segment_0;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire             p1_cpu_1_instruction_master_latency_counter;
  wire    [ 15: 0] p1_dbs_16_reg_segment_0;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_1_instruction_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  wire             r_3;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module | ~cpu_1_instruction_master_requests_cpu_1_jtag_debug_module) & (cpu_1_instruction_master_granted_cpu_1_jtag_debug_module | ~cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module) & ((~cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module | ~cpu_1_instruction_master_read | (1 & ~d1_cpu_1_jtag_debug_module_end_xfer & cpu_1_instruction_master_read)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_1_instruction_master_run = r_0 & r_1 & r_2 & r_3;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_1_instruction_master_qualified_request_nios_system_clock_0_in | ~cpu_1_instruction_master_requests_nios_system_clock_0_in) & ((~cpu_1_instruction_master_qualified_request_nios_system_clock_0_in | ~cpu_1_instruction_master_read | (1 & ~nios_system_clock_0_in_waitrequest_from_sa & (cpu_1_instruction_master_dbs_address[1]) & cpu_1_instruction_master_read)));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1 | ~cpu_1_instruction_master_requests_onchip_memory2_0_s1) & (cpu_1_instruction_master_granted_onchip_memory2_0_s1 | ~cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1) & ((~cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_1_instruction_master_read) | (1 & (cpu_1_instruction_master_read)))) & 1 & (cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1 | ~cpu_1_instruction_master_requests_onchip_memory2_1_s1) & (cpu_1_instruction_master_granted_onchip_memory2_1_s1 | ~cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1) & ((~cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_1_instruction_master_read) | (1 & (cpu_1_instruction_master_read)))) & 1 & (cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1 | ~cpu_1_instruction_master_requests_onchip_memory2_2_s1) & (cpu_1_instruction_master_granted_onchip_memory2_2_s1 | ~cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1) & ((~cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_1_instruction_master_read) | (1 & (cpu_1_instruction_master_read))));

  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1 | ~cpu_1_instruction_master_requests_onchip_memory2_3_s1) & (cpu_1_instruction_master_granted_onchip_memory2_3_s1 | ~cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1) & ((~cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_1_instruction_master_read) | (1 & (cpu_1_instruction_master_read)))) & 1 & (cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_1_instruction_master_requests_sram_0_avalon_sram_slave) & (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave | ~cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave) & ((~cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_1_instruction_master_read | (1 & (cpu_1_instruction_master_dbs_address[1]) & cpu_1_instruction_master_read)));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_1_instruction_master_address_to_slave = cpu_1_instruction_master_address[24 : 0];

  //cpu_1_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_1_instruction_master_read_but_no_slave_selected <= cpu_1_instruction_master_read & cpu_1_instruction_master_run & ~cpu_1_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_1_instruction_master_is_granted_some_slave = cpu_1_instruction_master_granted_cpu_1_jtag_debug_module |
    cpu_1_instruction_master_granted_nios_system_clock_0_in |
    cpu_1_instruction_master_granted_onchip_memory2_0_s1 |
    cpu_1_instruction_master_granted_onchip_memory2_1_s1 |
    cpu_1_instruction_master_granted_onchip_memory2_2_s1 |
    cpu_1_instruction_master_granted_onchip_memory2_3_s1 |
    cpu_1_instruction_master_granted_sram_0_avalon_sram_slave;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_1_instruction_master_readdatavalid = cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1 |
    cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1 |
    cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1 |
    cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1 |
    (cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave & dbs_rdv_counter_overflow);

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_1_instruction_master_readdatavalid = cpu_1_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_1_instruction_master_readdatavalid |
    cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module |
    cpu_1_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_1_instruction_master_readdatavalid |
    (cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in & dbs_counter_overflow) |
    cpu_1_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_1_instruction_master_readdatavalid |
    cpu_1_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_1_instruction_master_readdatavalid |
    cpu_1_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_1_instruction_master_readdatavalid |
    cpu_1_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_1_instruction_master_readdatavalid |
    cpu_1_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_1_instruction_master_readdatavalid;

  //cpu_1/instruction_master readdata mux, which is an e_mux
  assign cpu_1_instruction_master_readdata = ({32 {~(cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module & cpu_1_instruction_master_read)}} | cpu_1_jtag_debug_module_readdata_from_sa) &
    ({32 {~(cpu_1_instruction_master_qualified_request_nios_system_clock_0_in & cpu_1_instruction_master_read)}} | {nios_system_clock_0_in_readdata_from_sa[15 : 0],
    dbs_16_reg_segment_0}) &
    ({32 {~cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1}} | onchip_memory2_0_s1_readdata_from_sa) &
    ({32 {~cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1}} | onchip_memory2_1_s1_readdata_from_sa) &
    ({32 {~cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1}} | onchip_memory2_2_s1_readdata_from_sa) &
    ({32 {~cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1}} | onchip_memory2_3_s1_readdata_from_sa) &
    ({32 {~cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave}} | {sram_0_avalon_sram_slave_readdata_from_sa[15 : 0],
    dbs_latent_16_reg_segment_0});

  //actual waitrequest port, which is an e_assign
  assign cpu_1_instruction_master_waitrequest = ~cpu_1_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_instruction_master_latency_counter <= 0;
      else 
        cpu_1_instruction_master_latency_counter <= p1_cpu_1_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_1_instruction_master_latency_counter = ((cpu_1_instruction_master_run & cpu_1_instruction_master_read))? latency_load_value :
    (cpu_1_instruction_master_latency_counter)? cpu_1_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({1 {cpu_1_instruction_master_requests_onchip_memory2_0_s1}} & 1) |
    ({1 {cpu_1_instruction_master_requests_onchip_memory2_1_s1}} & 1) |
    ({1 {cpu_1_instruction_master_requests_onchip_memory2_2_s1}} & 1) |
    ({1 {cpu_1_instruction_master_requests_onchip_memory2_3_s1}} & 1);

  //input to dbs-16 stored 0, which is an e_mux
  assign p1_dbs_16_reg_segment_0 = nios_system_clock_0_in_readdata_from_sa;

  //dbs register for dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_16_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_1_instruction_master_dbs_address[1]) == 0))
          dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
    end


  //dbs count increment, which is an e_mux
  assign cpu_1_instruction_master_dbs_increment = (cpu_1_instruction_master_requests_nios_system_clock_0_in)? 2 :
    (cpu_1_instruction_master_requests_sram_0_avalon_sram_slave)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_1_instruction_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_1_instruction_master_dbs_address + cpu_1_instruction_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_instruction_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_1_instruction_master_dbs_address <= next_dbs_address;
    end


  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (cpu_1_instruction_master_granted_nios_system_clock_0_in & cpu_1_instruction_master_read & 1 & 1 & ~nios_system_clock_0_in_waitrequest_from_sa) |
    (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave & cpu_1_instruction_master_read & 1 & 1);

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = sram_0_avalon_sram_slave_readdata_from_sa;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_1_instruction_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_1_instruction_master_next_dbs_rdv_counter = cpu_1_instruction_master_dbs_rdv_counter + cpu_1_instruction_master_dbs_rdv_counter_inc;

  //cpu_1_instruction_master_rdv_inc_mux, which is an e_mux
  assign cpu_1_instruction_master_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_instruction_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_1_instruction_master_dbs_rdv_counter <= cpu_1_instruction_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_1_instruction_master_dbs_rdv_counter[1] & ~cpu_1_instruction_master_next_dbs_rdv_counter[1];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_1_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_instruction_master_address_last_time <= 0;
      else 
        cpu_1_instruction_master_address_last_time <= cpu_1_instruction_master_address;
    end


  //cpu_1/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_1_instruction_master_waitrequest & (cpu_1_instruction_master_read);
    end


  //cpu_1_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_1_instruction_master_address != cpu_1_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_1_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_1_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_instruction_master_read_last_time <= 0;
      else 
        cpu_1_instruction_master_read_last_time <= cpu_1_instruction_master_read;
    end


  //cpu_1_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_1_instruction_master_read != cpu_1_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_1_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_1_altera_nios_custom_instr_floating_point_inst_s1_arbitrator (
                                                                          // inputs:
                                                                           clk,
                                                                           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done,
                                                                           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result,
                                                                           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select,
                                                                           cpu_1_custom_instruction_master_multi_clk_en,
                                                                           cpu_1_custom_instruction_master_multi_dataa,
                                                                           cpu_1_custom_instruction_master_multi_datab,
                                                                           cpu_1_custom_instruction_master_multi_n,
                                                                           cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1,
                                                                           reset_n,

                                                                          // outputs:
                                                                           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_clk_en,
                                                                           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_dataa,
                                                                           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_datab,
                                                                           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa,
                                                                           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_n,
                                                                           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_reset,
                                                                           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa,
                                                                           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_start
                                                                        )
;

  output           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  output  [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  output  [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_datab;
  output           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  output  [  1: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_n;
  output           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_reset;
  output  [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  output           cpu_1_altera_nios_custom_instr_floating_point_inst_s1_start;
  input            clk;
  input            cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done;
  input   [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result;
  input            cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select;
  input            cpu_1_custom_instruction_master_multi_clk_en;
  input   [ 31: 0] cpu_1_custom_instruction_master_multi_dataa;
  input   [ 31: 0] cpu_1_custom_instruction_master_multi_datab;
  input   [  7: 0] cpu_1_custom_instruction_master_multi_n;
  input            cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1;
  input            reset_n;

  wire             cpu_1_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  wire    [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  wire    [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_datab;
  wire             cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  wire    [  1: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_n;
  wire             cpu_1_altera_nios_custom_instr_floating_point_inst_s1_reset;
  wire    [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  wire             cpu_1_altera_nios_custom_instr_floating_point_inst_s1_start;
  assign cpu_1_altera_nios_custom_instr_floating_point_inst_s1_clk_en = cpu_1_custom_instruction_master_multi_clk_en;
  assign cpu_1_altera_nios_custom_instr_floating_point_inst_s1_dataa = cpu_1_custom_instruction_master_multi_dataa;
  assign cpu_1_altera_nios_custom_instr_floating_point_inst_s1_datab = cpu_1_custom_instruction_master_multi_datab;
  assign cpu_1_altera_nios_custom_instr_floating_point_inst_s1_n = cpu_1_custom_instruction_master_multi_n;
  assign cpu_1_altera_nios_custom_instr_floating_point_inst_s1_start = cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1;
  //assign cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa = cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa = cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result;

  //assign cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa = cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa = cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done;

  //cpu_1_altera_nios_custom_instr_floating_point_inst/s1 local reset_n, which is an e_assign
  assign cpu_1_altera_nios_custom_instr_floating_point_inst_s1_reset = ~reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_2_jtag_debug_module_arbitrator (
                                            // inputs:
                                             clk,
                                             cpu_2_data_master_address_to_slave,
                                             cpu_2_data_master_byteenable,
                                             cpu_2_data_master_debugaccess,
                                             cpu_2_data_master_latency_counter,
                                             cpu_2_data_master_read,
                                             cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                             cpu_2_data_master_write,
                                             cpu_2_data_master_writedata,
                                             cpu_2_instruction_master_address_to_slave,
                                             cpu_2_instruction_master_latency_counter,
                                             cpu_2_instruction_master_read,
                                             cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                             cpu_2_jtag_debug_module_readdata,
                                             cpu_2_jtag_debug_module_resetrequest,
                                             reset_n,

                                            // outputs:
                                             cpu_2_data_master_granted_cpu_2_jtag_debug_module,
                                             cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module,
                                             cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module,
                                             cpu_2_data_master_requests_cpu_2_jtag_debug_module,
                                             cpu_2_instruction_master_granted_cpu_2_jtag_debug_module,
                                             cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module,
                                             cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module,
                                             cpu_2_instruction_master_requests_cpu_2_jtag_debug_module,
                                             cpu_2_jtag_debug_module_address,
                                             cpu_2_jtag_debug_module_begintransfer,
                                             cpu_2_jtag_debug_module_byteenable,
                                             cpu_2_jtag_debug_module_chipselect,
                                             cpu_2_jtag_debug_module_debugaccess,
                                             cpu_2_jtag_debug_module_readdata_from_sa,
                                             cpu_2_jtag_debug_module_resetrequest_from_sa,
                                             cpu_2_jtag_debug_module_write,
                                             cpu_2_jtag_debug_module_writedata,
                                             d1_cpu_2_jtag_debug_module_end_xfer
                                          )
;

  output           cpu_2_data_master_granted_cpu_2_jtag_debug_module;
  output           cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module;
  output           cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module;
  output           cpu_2_data_master_requests_cpu_2_jtag_debug_module;
  output           cpu_2_instruction_master_granted_cpu_2_jtag_debug_module;
  output           cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module;
  output           cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module;
  output           cpu_2_instruction_master_requests_cpu_2_jtag_debug_module;
  output  [  8: 0] cpu_2_jtag_debug_module_address;
  output           cpu_2_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_2_jtag_debug_module_byteenable;
  output           cpu_2_jtag_debug_module_chipselect;
  output           cpu_2_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_2_jtag_debug_module_readdata_from_sa;
  output           cpu_2_jtag_debug_module_resetrequest_from_sa;
  output           cpu_2_jtag_debug_module_write;
  output  [ 31: 0] cpu_2_jtag_debug_module_writedata;
  output           d1_cpu_2_jtag_debug_module_end_xfer;
  input            clk;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input   [  3: 0] cpu_2_data_master_byteenable;
  input            cpu_2_data_master_debugaccess;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_2_instruction_master_address_to_slave;
  input            cpu_2_instruction_master_latency_counter;
  input            cpu_2_instruction_master_read;
  input            cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 31: 0] cpu_2_jtag_debug_module_readdata;
  input            cpu_2_jtag_debug_module_resetrequest;
  input            reset_n;

  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_cpu_2_jtag_debug_module;
  wire             cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module;
  wire             cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module;
  wire             cpu_2_data_master_requests_cpu_2_jtag_debug_module;
  wire             cpu_2_data_master_saved_grant_cpu_2_jtag_debug_module;
  wire             cpu_2_instruction_master_arbiterlock;
  wire             cpu_2_instruction_master_arbiterlock2;
  wire             cpu_2_instruction_master_continuerequest;
  wire             cpu_2_instruction_master_granted_cpu_2_jtag_debug_module;
  wire             cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module;
  wire             cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module;
  wire             cpu_2_instruction_master_requests_cpu_2_jtag_debug_module;
  wire             cpu_2_instruction_master_saved_grant_cpu_2_jtag_debug_module;
  wire    [  8: 0] cpu_2_jtag_debug_module_address;
  wire             cpu_2_jtag_debug_module_allgrants;
  wire             cpu_2_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_2_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_2_jtag_debug_module_any_continuerequest;
  reg     [  1: 0] cpu_2_jtag_debug_module_arb_addend;
  wire             cpu_2_jtag_debug_module_arb_counter_enable;
  reg     [  2: 0] cpu_2_jtag_debug_module_arb_share_counter;
  wire    [  2: 0] cpu_2_jtag_debug_module_arb_share_counter_next_value;
  wire    [  2: 0] cpu_2_jtag_debug_module_arb_share_set_values;
  wire    [  1: 0] cpu_2_jtag_debug_module_arb_winner;
  wire             cpu_2_jtag_debug_module_arbitration_holdoff_internal;
  wire             cpu_2_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_2_jtag_debug_module_begins_xfer;
  wire             cpu_2_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_2_jtag_debug_module_byteenable;
  wire             cpu_2_jtag_debug_module_chipselect;
  wire    [  3: 0] cpu_2_jtag_debug_module_chosen_master_double_vector;
  wire    [  1: 0] cpu_2_jtag_debug_module_chosen_master_rot_left;
  wire             cpu_2_jtag_debug_module_debugaccess;
  wire             cpu_2_jtag_debug_module_end_xfer;
  wire             cpu_2_jtag_debug_module_firsttransfer;
  wire    [  1: 0] cpu_2_jtag_debug_module_grant_vector;
  wire             cpu_2_jtag_debug_module_in_a_read_cycle;
  wire             cpu_2_jtag_debug_module_in_a_write_cycle;
  wire    [  1: 0] cpu_2_jtag_debug_module_master_qreq_vector;
  wire             cpu_2_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_2_jtag_debug_module_readdata_from_sa;
  reg              cpu_2_jtag_debug_module_reg_firsttransfer;
  wire             cpu_2_jtag_debug_module_resetrequest_from_sa;
  reg     [  1: 0] cpu_2_jtag_debug_module_saved_chosen_master_vector;
  reg              cpu_2_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_2_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_2_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_2_jtag_debug_module_waits_for_read;
  wire             cpu_2_jtag_debug_module_waits_for_write;
  wire             cpu_2_jtag_debug_module_write;
  wire    [ 31: 0] cpu_2_jtag_debug_module_writedata;
  reg              d1_cpu_2_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_2_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_2_data_master_granted_slave_cpu_2_jtag_debug_module;
  reg              last_cycle_cpu_2_instruction_master_granted_slave_cpu_2_jtag_debug_module;
  wire    [ 24: 0] shifted_address_to_cpu_2_jtag_debug_module_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_cpu_2_jtag_debug_module_from_cpu_2_instruction_master;
  wire             wait_for_cpu_2_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_2_jtag_debug_module_end_xfer;
    end


  assign cpu_2_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module | cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module));
  //assign cpu_2_jtag_debug_module_readdata_from_sa = cpu_2_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_2_jtag_debug_module_readdata_from_sa = cpu_2_jtag_debug_module_readdata;

  assign cpu_2_data_master_requests_cpu_2_jtag_debug_module = ({cpu_2_data_master_address_to_slave[24 : 11] , 11'b0} == 25'h1800) & (cpu_2_data_master_read | cpu_2_data_master_write);
  //cpu_2_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_2_jtag_debug_module_arb_share_set_values = 1;

  //cpu_2_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_2_jtag_debug_module_non_bursting_master_requests = cpu_2_data_master_requests_cpu_2_jtag_debug_module |
    cpu_2_instruction_master_requests_cpu_2_jtag_debug_module |
    cpu_2_data_master_requests_cpu_2_jtag_debug_module |
    cpu_2_instruction_master_requests_cpu_2_jtag_debug_module;

  //cpu_2_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_2_jtag_debug_module_any_bursting_master_saved_grant = 0;

  //cpu_2_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_2_jtag_debug_module_arb_share_counter_next_value = cpu_2_jtag_debug_module_firsttransfer ? (cpu_2_jtag_debug_module_arb_share_set_values - 1) : |cpu_2_jtag_debug_module_arb_share_counter ? (cpu_2_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_2_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_2_jtag_debug_module_allgrants = (|cpu_2_jtag_debug_module_grant_vector) |
    (|cpu_2_jtag_debug_module_grant_vector) |
    (|cpu_2_jtag_debug_module_grant_vector) |
    (|cpu_2_jtag_debug_module_grant_vector);

  //cpu_2_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_2_jtag_debug_module_end_xfer = ~(cpu_2_jtag_debug_module_waits_for_read | cpu_2_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_2_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_2_jtag_debug_module = cpu_2_jtag_debug_module_end_xfer & (~cpu_2_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_2_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_2_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_2_jtag_debug_module & cpu_2_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_2_jtag_debug_module & ~cpu_2_jtag_debug_module_non_bursting_master_requests);

  //cpu_2_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_2_jtag_debug_module_arb_counter_enable)
          cpu_2_jtag_debug_module_arb_share_counter <= cpu_2_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_2_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_2_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_2_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_2_jtag_debug_module & ~cpu_2_jtag_debug_module_non_bursting_master_requests))
          cpu_2_jtag_debug_module_slavearbiterlockenable <= |cpu_2_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_2/data_master cpu_2/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = cpu_2_jtag_debug_module_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_2_jtag_debug_module_slavearbiterlockenable2 = |cpu_2_jtag_debug_module_arb_share_counter_next_value;

  //cpu_2/data_master cpu_2/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = cpu_2_jtag_debug_module_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/instruction_master cpu_2/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock = cpu_2_jtag_debug_module_slavearbiterlockenable & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master cpu_2/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock2 = cpu_2_jtag_debug_module_slavearbiterlockenable2 & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master granted cpu_2/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_instruction_master_granted_slave_cpu_2_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_2_instruction_master_granted_slave_cpu_2_jtag_debug_module <= cpu_2_instruction_master_saved_grant_cpu_2_jtag_debug_module ? 1 : (cpu_2_jtag_debug_module_arbitration_holdoff_internal | ~cpu_2_instruction_master_requests_cpu_2_jtag_debug_module) ? 0 : last_cycle_cpu_2_instruction_master_granted_slave_cpu_2_jtag_debug_module;
    end


  //cpu_2_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_2_instruction_master_continuerequest = last_cycle_cpu_2_instruction_master_granted_slave_cpu_2_jtag_debug_module & cpu_2_instruction_master_requests_cpu_2_jtag_debug_module;

  //cpu_2_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_2_jtag_debug_module_any_continuerequest = cpu_2_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest;

  assign cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module = cpu_2_data_master_requests_cpu_2_jtag_debug_module & ~((cpu_2_data_master_read & ((cpu_2_data_master_latency_counter != 0) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_2_instruction_master_arbiterlock);
  //local readdatavalid cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module, which is an e_mux
  assign cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module = cpu_2_data_master_granted_cpu_2_jtag_debug_module & cpu_2_data_master_read & ~cpu_2_jtag_debug_module_waits_for_read;

  //cpu_2_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_2_jtag_debug_module_writedata = cpu_2_data_master_writedata;

  assign cpu_2_instruction_master_requests_cpu_2_jtag_debug_module = (({cpu_2_instruction_master_address_to_slave[24 : 11] , 11'b0} == 25'h1800) & (cpu_2_instruction_master_read)) & cpu_2_instruction_master_read;
  //cpu_2/data_master granted cpu_2/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_cpu_2_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_cpu_2_jtag_debug_module <= cpu_2_data_master_saved_grant_cpu_2_jtag_debug_module ? 1 : (cpu_2_jtag_debug_module_arbitration_holdoff_internal | ~cpu_2_data_master_requests_cpu_2_jtag_debug_module) ? 0 : last_cycle_cpu_2_data_master_granted_slave_cpu_2_jtag_debug_module;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = last_cycle_cpu_2_data_master_granted_slave_cpu_2_jtag_debug_module & cpu_2_data_master_requests_cpu_2_jtag_debug_module;

  assign cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module = cpu_2_instruction_master_requests_cpu_2_jtag_debug_module & ~((cpu_2_instruction_master_read & ((cpu_2_instruction_master_latency_counter != 0) | (|cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_2_data_master_arbiterlock);
  //local readdatavalid cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module, which is an e_mux
  assign cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module = cpu_2_instruction_master_granted_cpu_2_jtag_debug_module & cpu_2_instruction_master_read & ~cpu_2_jtag_debug_module_waits_for_read;

  //allow new arb cycle for cpu_2/jtag_debug_module, which is an e_assign
  assign cpu_2_jtag_debug_module_allow_new_arb_cycle = ~cpu_2_data_master_arbiterlock & ~cpu_2_instruction_master_arbiterlock;

  //cpu_2/instruction_master assignment into master qualified-requests vector for cpu_2/jtag_debug_module, which is an e_assign
  assign cpu_2_jtag_debug_module_master_qreq_vector[0] = cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module;

  //cpu_2/instruction_master grant cpu_2/jtag_debug_module, which is an e_assign
  assign cpu_2_instruction_master_granted_cpu_2_jtag_debug_module = cpu_2_jtag_debug_module_grant_vector[0];

  //cpu_2/instruction_master saved-grant cpu_2/jtag_debug_module, which is an e_assign
  assign cpu_2_instruction_master_saved_grant_cpu_2_jtag_debug_module = cpu_2_jtag_debug_module_arb_winner[0] && cpu_2_instruction_master_requests_cpu_2_jtag_debug_module;

  //cpu_2/data_master assignment into master qualified-requests vector for cpu_2/jtag_debug_module, which is an e_assign
  assign cpu_2_jtag_debug_module_master_qreq_vector[1] = cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module;

  //cpu_2/data_master grant cpu_2/jtag_debug_module, which is an e_assign
  assign cpu_2_data_master_granted_cpu_2_jtag_debug_module = cpu_2_jtag_debug_module_grant_vector[1];

  //cpu_2/data_master saved-grant cpu_2/jtag_debug_module, which is an e_assign
  assign cpu_2_data_master_saved_grant_cpu_2_jtag_debug_module = cpu_2_jtag_debug_module_arb_winner[1] && cpu_2_data_master_requests_cpu_2_jtag_debug_module;

  //cpu_2/jtag_debug_module chosen-master double-vector, which is an e_assign
  assign cpu_2_jtag_debug_module_chosen_master_double_vector = {cpu_2_jtag_debug_module_master_qreq_vector, cpu_2_jtag_debug_module_master_qreq_vector} & ({~cpu_2_jtag_debug_module_master_qreq_vector, ~cpu_2_jtag_debug_module_master_qreq_vector} + cpu_2_jtag_debug_module_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_2_jtag_debug_module_arb_winner = (cpu_2_jtag_debug_module_allow_new_arb_cycle & | cpu_2_jtag_debug_module_grant_vector) ? cpu_2_jtag_debug_module_grant_vector : cpu_2_jtag_debug_module_saved_chosen_master_vector;

  //saved cpu_2_jtag_debug_module_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_jtag_debug_module_saved_chosen_master_vector <= 0;
      else if (cpu_2_jtag_debug_module_allow_new_arb_cycle)
          cpu_2_jtag_debug_module_saved_chosen_master_vector <= |cpu_2_jtag_debug_module_grant_vector ? cpu_2_jtag_debug_module_grant_vector : cpu_2_jtag_debug_module_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_2_jtag_debug_module_grant_vector = {(cpu_2_jtag_debug_module_chosen_master_double_vector[1] | cpu_2_jtag_debug_module_chosen_master_double_vector[3]),
    (cpu_2_jtag_debug_module_chosen_master_double_vector[0] | cpu_2_jtag_debug_module_chosen_master_double_vector[2])};

  //cpu_2/jtag_debug_module chosen master rotated left, which is an e_assign
  assign cpu_2_jtag_debug_module_chosen_master_rot_left = (cpu_2_jtag_debug_module_arb_winner << 1) ? (cpu_2_jtag_debug_module_arb_winner << 1) : 1;

  //cpu_2/jtag_debug_module's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_jtag_debug_module_arb_addend <= 1;
      else if (|cpu_2_jtag_debug_module_grant_vector)
          cpu_2_jtag_debug_module_arb_addend <= cpu_2_jtag_debug_module_end_xfer? cpu_2_jtag_debug_module_chosen_master_rot_left : cpu_2_jtag_debug_module_grant_vector;
    end


  assign cpu_2_jtag_debug_module_begintransfer = cpu_2_jtag_debug_module_begins_xfer;
  //assign cpu_2_jtag_debug_module_resetrequest_from_sa = cpu_2_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_2_jtag_debug_module_resetrequest_from_sa = cpu_2_jtag_debug_module_resetrequest;

  assign cpu_2_jtag_debug_module_chipselect = cpu_2_data_master_granted_cpu_2_jtag_debug_module | cpu_2_instruction_master_granted_cpu_2_jtag_debug_module;
  //cpu_2_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_2_jtag_debug_module_firsttransfer = cpu_2_jtag_debug_module_begins_xfer ? cpu_2_jtag_debug_module_unreg_firsttransfer : cpu_2_jtag_debug_module_reg_firsttransfer;

  //cpu_2_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_2_jtag_debug_module_unreg_firsttransfer = ~(cpu_2_jtag_debug_module_slavearbiterlockenable & cpu_2_jtag_debug_module_any_continuerequest);

  //cpu_2_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_2_jtag_debug_module_begins_xfer)
          cpu_2_jtag_debug_module_reg_firsttransfer <= cpu_2_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_2_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_2_jtag_debug_module_beginbursttransfer_internal = cpu_2_jtag_debug_module_begins_xfer;

  //cpu_2_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_2_jtag_debug_module_arbitration_holdoff_internal = cpu_2_jtag_debug_module_begins_xfer & cpu_2_jtag_debug_module_firsttransfer;

  //cpu_2_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_2_jtag_debug_module_write = cpu_2_data_master_granted_cpu_2_jtag_debug_module & cpu_2_data_master_write;

  assign shifted_address_to_cpu_2_jtag_debug_module_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  //cpu_2_jtag_debug_module_address mux, which is an e_mux
  assign cpu_2_jtag_debug_module_address = (cpu_2_data_master_granted_cpu_2_jtag_debug_module)? (shifted_address_to_cpu_2_jtag_debug_module_from_cpu_2_data_master >> 2) :
    (shifted_address_to_cpu_2_jtag_debug_module_from_cpu_2_instruction_master >> 2);

  assign shifted_address_to_cpu_2_jtag_debug_module_from_cpu_2_instruction_master = cpu_2_instruction_master_address_to_slave;
  //d1_cpu_2_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_2_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_2_jtag_debug_module_end_xfer <= cpu_2_jtag_debug_module_end_xfer;
    end


  //cpu_2_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_2_jtag_debug_module_waits_for_read = cpu_2_jtag_debug_module_in_a_read_cycle & cpu_2_jtag_debug_module_begins_xfer;

  //cpu_2_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_2_jtag_debug_module_in_a_read_cycle = (cpu_2_data_master_granted_cpu_2_jtag_debug_module & cpu_2_data_master_read) | (cpu_2_instruction_master_granted_cpu_2_jtag_debug_module & cpu_2_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_2_jtag_debug_module_in_a_read_cycle;

  //cpu_2_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_2_jtag_debug_module_waits_for_write = cpu_2_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_2_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_2_jtag_debug_module_in_a_write_cycle = cpu_2_data_master_granted_cpu_2_jtag_debug_module & cpu_2_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_2_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_2_jtag_debug_module_counter = 0;
  //cpu_2_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_2_jtag_debug_module_byteenable = (cpu_2_data_master_granted_cpu_2_jtag_debug_module)? cpu_2_data_master_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_2_jtag_debug_module_debugaccess = (cpu_2_data_master_granted_cpu_2_jtag_debug_module)? cpu_2_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_2/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_2_data_master_granted_cpu_2_jtag_debug_module + cpu_2_instruction_master_granted_cpu_2_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_2_data_master_saved_grant_cpu_2_jtag_debug_module + cpu_2_instruction_master_saved_grant_cpu_2_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_2_custom_instruction_master_arbitrator (
                                                    // inputs:
                                                     clk,
                                                     cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa,
                                                     cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa,
                                                     cpu_2_custom_instruction_master_multi_start,
                                                     reset_n,

                                                    // outputs:
                                                     cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select,
                                                     cpu_2_custom_instruction_master_multi_done,
                                                     cpu_2_custom_instruction_master_multi_result,
                                                     cpu_2_custom_instruction_master_reset_n,
                                                     cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1
                                                  )
;

  output           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select;
  output           cpu_2_custom_instruction_master_multi_done;
  output  [ 31: 0] cpu_2_custom_instruction_master_multi_result;
  output           cpu_2_custom_instruction_master_reset_n;
  output           cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1;
  input            clk;
  input            cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  input   [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  input            cpu_2_custom_instruction_master_multi_start;
  input            reset_n;

  wire             cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select;
  wire             cpu_2_custom_instruction_master_multi_done;
  wire    [ 31: 0] cpu_2_custom_instruction_master_multi_result;
  wire             cpu_2_custom_instruction_master_reset_n;
  wire             cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1;
  assign cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select = 1'b1;
  assign cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1 = cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select & cpu_2_custom_instruction_master_multi_start;
  //cpu_2_custom_instruction_master_multi_result mux, which is an e_mux
  assign cpu_2_custom_instruction_master_multi_result = {32 {cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select}} & cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;

  //multi_done mux, which is an e_mux
  assign cpu_2_custom_instruction_master_multi_done = {1 {cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select}} & cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;

  //cpu_2_custom_instruction_master_reset_n local reset_n, which is an e_assign
  assign cpu_2_custom_instruction_master_reset_n = reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_2_data_master_arbitrator (
                                      // inputs:
                                       clk,
                                       cpu_2_data_master_address,
                                       cpu_2_data_master_byteenable,
                                       cpu_2_data_master_byteenable_nios_system_clock_10_in,
                                       cpu_2_data_master_byteenable_nios_system_clock_5_in,
                                       cpu_2_data_master_byteenable_sram_0_avalon_sram_slave,
                                       cpu_2_data_master_granted_cpu_2_jtag_debug_module,
                                       cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave,
                                       cpu_2_data_master_granted_keys_s1,
                                       cpu_2_data_master_granted_mailbox_0_s1,
                                       cpu_2_data_master_granted_mailbox_1_s1,
                                       cpu_2_data_master_granted_mailbox_2_s1,
                                       cpu_2_data_master_granted_mailbox_3_s1,
                                       cpu_2_data_master_granted_nios_system_clock_10_in,
                                       cpu_2_data_master_granted_nios_system_clock_5_in,
                                       cpu_2_data_master_granted_onchip_memory2_0_s1,
                                       cpu_2_data_master_granted_onchip_memory2_1_s1,
                                       cpu_2_data_master_granted_onchip_memory2_2_s1,
                                       cpu_2_data_master_granted_onchip_memory2_3_s1,
                                       cpu_2_data_master_granted_performance_counter_0_control_slave,
                                       cpu_2_data_master_granted_sram_0_avalon_sram_slave,
                                       cpu_2_data_master_granted_sysid_control_slave,
                                       cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module,
                                       cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave,
                                       cpu_2_data_master_qualified_request_keys_s1,
                                       cpu_2_data_master_qualified_request_mailbox_0_s1,
                                       cpu_2_data_master_qualified_request_mailbox_1_s1,
                                       cpu_2_data_master_qualified_request_mailbox_2_s1,
                                       cpu_2_data_master_qualified_request_mailbox_3_s1,
                                       cpu_2_data_master_qualified_request_nios_system_clock_10_in,
                                       cpu_2_data_master_qualified_request_nios_system_clock_5_in,
                                       cpu_2_data_master_qualified_request_onchip_memory2_0_s1,
                                       cpu_2_data_master_qualified_request_onchip_memory2_1_s1,
                                       cpu_2_data_master_qualified_request_onchip_memory2_2_s1,
                                       cpu_2_data_master_qualified_request_onchip_memory2_3_s1,
                                       cpu_2_data_master_qualified_request_performance_counter_0_control_slave,
                                       cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave,
                                       cpu_2_data_master_qualified_request_sysid_control_slave,
                                       cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_2_data_master_read,
                                       cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module,
                                       cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave,
                                       cpu_2_data_master_read_data_valid_keys_s1,
                                       cpu_2_data_master_read_data_valid_mailbox_0_s1,
                                       cpu_2_data_master_read_data_valid_mailbox_1_s1,
                                       cpu_2_data_master_read_data_valid_mailbox_2_s1,
                                       cpu_2_data_master_read_data_valid_mailbox_3_s1,
                                       cpu_2_data_master_read_data_valid_nios_system_clock_10_in,
                                       cpu_2_data_master_read_data_valid_nios_system_clock_5_in,
                                       cpu_2_data_master_read_data_valid_onchip_memory2_0_s1,
                                       cpu_2_data_master_read_data_valid_onchip_memory2_1_s1,
                                       cpu_2_data_master_read_data_valid_onchip_memory2_2_s1,
                                       cpu_2_data_master_read_data_valid_onchip_memory2_3_s1,
                                       cpu_2_data_master_read_data_valid_performance_counter_0_control_slave,
                                       cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave,
                                       cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                       cpu_2_data_master_read_data_valid_sysid_control_slave,
                                       cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_2_data_master_requests_cpu_2_jtag_debug_module,
                                       cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave,
                                       cpu_2_data_master_requests_keys_s1,
                                       cpu_2_data_master_requests_mailbox_0_s1,
                                       cpu_2_data_master_requests_mailbox_1_s1,
                                       cpu_2_data_master_requests_mailbox_2_s1,
                                       cpu_2_data_master_requests_mailbox_3_s1,
                                       cpu_2_data_master_requests_nios_system_clock_10_in,
                                       cpu_2_data_master_requests_nios_system_clock_5_in,
                                       cpu_2_data_master_requests_onchip_memory2_0_s1,
                                       cpu_2_data_master_requests_onchip_memory2_1_s1,
                                       cpu_2_data_master_requests_onchip_memory2_2_s1,
                                       cpu_2_data_master_requests_onchip_memory2_3_s1,
                                       cpu_2_data_master_requests_performance_counter_0_control_slave,
                                       cpu_2_data_master_requests_sram_0_avalon_sram_slave,
                                       cpu_2_data_master_requests_sysid_control_slave,
                                       cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_2_data_master_write,
                                       cpu_2_data_master_writedata,
                                       cpu_2_jtag_debug_module_readdata_from_sa,
                                       d1_cpu_2_jtag_debug_module_end_xfer,
                                       d1_jtag_uart_2_avalon_jtag_slave_end_xfer,
                                       d1_keys_s1_end_xfer,
                                       d1_mailbox_0_s1_end_xfer,
                                       d1_mailbox_1_s1_end_xfer,
                                       d1_mailbox_2_s1_end_xfer,
                                       d1_mailbox_3_s1_end_xfer,
                                       d1_nios_system_clock_10_in_end_xfer,
                                       d1_nios_system_clock_5_in_end_xfer,
                                       d1_onchip_memory2_0_s1_end_xfer,
                                       d1_onchip_memory2_1_s1_end_xfer,
                                       d1_onchip_memory2_2_s1_end_xfer,
                                       d1_onchip_memory2_3_s1_end_xfer,
                                       d1_performance_counter_0_control_slave_end_xfer,
                                       d1_sram_0_avalon_sram_slave_end_xfer,
                                       d1_sysid_control_slave_end_xfer,
                                       d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer,
                                       jtag_uart_2_avalon_jtag_slave_irq_from_sa,
                                       jtag_uart_2_avalon_jtag_slave_readdata_from_sa,
                                       jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa,
                                       keys_s1_readdata_from_sa,
                                       mailbox_0_s1_readdata_from_sa,
                                       mailbox_1_s1_readdata_from_sa,
                                       mailbox_2_s1_readdata_from_sa,
                                       mailbox_3_s1_readdata_from_sa,
                                       nios_system_clock_10_in_readdata_from_sa,
                                       nios_system_clock_10_in_waitrequest_from_sa,
                                       nios_system_clock_5_in_readdata_from_sa,
                                       nios_system_clock_5_in_waitrequest_from_sa,
                                       onchip_memory2_0_s1_readdata_from_sa,
                                       onchip_memory2_1_s1_readdata_from_sa,
                                       onchip_memory2_2_s1_readdata_from_sa,
                                       onchip_memory2_3_s1_readdata_from_sa,
                                       performance_counter_0_control_slave_readdata_from_sa,
                                       reset_n,
                                       sram_0_avalon_sram_slave_readdata_from_sa,
                                       sysid_control_slave_readdata_from_sa,
                                       video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa,

                                      // outputs:
                                       cpu_2_data_master_address_to_slave,
                                       cpu_2_data_master_dbs_address,
                                       cpu_2_data_master_dbs_write_16,
                                       cpu_2_data_master_dbs_write_8,
                                       cpu_2_data_master_irq,
                                       cpu_2_data_master_latency_counter,
                                       cpu_2_data_master_readdata,
                                       cpu_2_data_master_readdatavalid,
                                       cpu_2_data_master_waitrequest
                                    )
;

  output  [ 24: 0] cpu_2_data_master_address_to_slave;
  output  [  1: 0] cpu_2_data_master_dbs_address;
  output  [ 15: 0] cpu_2_data_master_dbs_write_16;
  output  [  7: 0] cpu_2_data_master_dbs_write_8;
  output  [ 31: 0] cpu_2_data_master_irq;
  output           cpu_2_data_master_latency_counter;
  output  [ 31: 0] cpu_2_data_master_readdata;
  output           cpu_2_data_master_readdatavalid;
  output           cpu_2_data_master_waitrequest;
  input            clk;
  input   [ 24: 0] cpu_2_data_master_address;
  input   [  3: 0] cpu_2_data_master_byteenable;
  input            cpu_2_data_master_byteenable_nios_system_clock_10_in;
  input   [  1: 0] cpu_2_data_master_byteenable_nios_system_clock_5_in;
  input   [  1: 0] cpu_2_data_master_byteenable_sram_0_avalon_sram_slave;
  input            cpu_2_data_master_granted_cpu_2_jtag_debug_module;
  input            cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave;
  input            cpu_2_data_master_granted_keys_s1;
  input            cpu_2_data_master_granted_mailbox_0_s1;
  input            cpu_2_data_master_granted_mailbox_1_s1;
  input            cpu_2_data_master_granted_mailbox_2_s1;
  input            cpu_2_data_master_granted_mailbox_3_s1;
  input            cpu_2_data_master_granted_nios_system_clock_10_in;
  input            cpu_2_data_master_granted_nios_system_clock_5_in;
  input            cpu_2_data_master_granted_onchip_memory2_0_s1;
  input            cpu_2_data_master_granted_onchip_memory2_1_s1;
  input            cpu_2_data_master_granted_onchip_memory2_2_s1;
  input            cpu_2_data_master_granted_onchip_memory2_3_s1;
  input            cpu_2_data_master_granted_performance_counter_0_control_slave;
  input            cpu_2_data_master_granted_sram_0_avalon_sram_slave;
  input            cpu_2_data_master_granted_sysid_control_slave;
  input            cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module;
  input            cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave;
  input            cpu_2_data_master_qualified_request_keys_s1;
  input            cpu_2_data_master_qualified_request_mailbox_0_s1;
  input            cpu_2_data_master_qualified_request_mailbox_1_s1;
  input            cpu_2_data_master_qualified_request_mailbox_2_s1;
  input            cpu_2_data_master_qualified_request_mailbox_3_s1;
  input            cpu_2_data_master_qualified_request_nios_system_clock_10_in;
  input            cpu_2_data_master_qualified_request_nios_system_clock_5_in;
  input            cpu_2_data_master_qualified_request_onchip_memory2_0_s1;
  input            cpu_2_data_master_qualified_request_onchip_memory2_1_s1;
  input            cpu_2_data_master_qualified_request_onchip_memory2_2_s1;
  input            cpu_2_data_master_qualified_request_onchip_memory2_3_s1;
  input            cpu_2_data_master_qualified_request_performance_counter_0_control_slave;
  input            cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave;
  input            cpu_2_data_master_qualified_request_sysid_control_slave;
  input            cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module;
  input            cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave;
  input            cpu_2_data_master_read_data_valid_keys_s1;
  input            cpu_2_data_master_read_data_valid_mailbox_0_s1;
  input            cpu_2_data_master_read_data_valid_mailbox_1_s1;
  input            cpu_2_data_master_read_data_valid_mailbox_2_s1;
  input            cpu_2_data_master_read_data_valid_mailbox_3_s1;
  input            cpu_2_data_master_read_data_valid_nios_system_clock_10_in;
  input            cpu_2_data_master_read_data_valid_nios_system_clock_5_in;
  input            cpu_2_data_master_read_data_valid_onchip_memory2_0_s1;
  input            cpu_2_data_master_read_data_valid_onchip_memory2_1_s1;
  input            cpu_2_data_master_read_data_valid_onchip_memory2_2_s1;
  input            cpu_2_data_master_read_data_valid_onchip_memory2_3_s1;
  input            cpu_2_data_master_read_data_valid_performance_counter_0_control_slave;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_read_data_valid_sysid_control_slave;
  input            cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_2_data_master_requests_cpu_2_jtag_debug_module;
  input            cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave;
  input            cpu_2_data_master_requests_keys_s1;
  input            cpu_2_data_master_requests_mailbox_0_s1;
  input            cpu_2_data_master_requests_mailbox_1_s1;
  input            cpu_2_data_master_requests_mailbox_2_s1;
  input            cpu_2_data_master_requests_mailbox_3_s1;
  input            cpu_2_data_master_requests_nios_system_clock_10_in;
  input            cpu_2_data_master_requests_nios_system_clock_5_in;
  input            cpu_2_data_master_requests_onchip_memory2_0_s1;
  input            cpu_2_data_master_requests_onchip_memory2_1_s1;
  input            cpu_2_data_master_requests_onchip_memory2_2_s1;
  input            cpu_2_data_master_requests_onchip_memory2_3_s1;
  input            cpu_2_data_master_requests_performance_counter_0_control_slave;
  input            cpu_2_data_master_requests_sram_0_avalon_sram_slave;
  input            cpu_2_data_master_requests_sysid_control_slave;
  input            cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 31: 0] cpu_2_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_2_jtag_debug_module_end_xfer;
  input            d1_jtag_uart_2_avalon_jtag_slave_end_xfer;
  input            d1_keys_s1_end_xfer;
  input            d1_mailbox_0_s1_end_xfer;
  input            d1_mailbox_1_s1_end_xfer;
  input            d1_mailbox_2_s1_end_xfer;
  input            d1_mailbox_3_s1_end_xfer;
  input            d1_nios_system_clock_10_in_end_xfer;
  input            d1_nios_system_clock_5_in_end_xfer;
  input            d1_onchip_memory2_0_s1_end_xfer;
  input            d1_onchip_memory2_1_s1_end_xfer;
  input            d1_onchip_memory2_2_s1_end_xfer;
  input            d1_onchip_memory2_3_s1_end_xfer;
  input            d1_performance_counter_0_control_slave_end_xfer;
  input            d1_sram_0_avalon_sram_slave_end_xfer;
  input            d1_sysid_control_slave_end_xfer;
  input            d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer;
  input            jtag_uart_2_avalon_jtag_slave_irq_from_sa;
  input   [ 31: 0] jtag_uart_2_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa;
  input   [ 31: 0] keys_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_0_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_1_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_2_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_3_s1_readdata_from_sa;
  input   [  7: 0] nios_system_clock_10_in_readdata_from_sa;
  input            nios_system_clock_10_in_waitrequest_from_sa;
  input   [ 15: 0] nios_system_clock_5_in_readdata_from_sa;
  input            nios_system_clock_5_in_waitrequest_from_sa;
  input   [ 31: 0] onchip_memory2_0_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_1_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_2_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_3_s1_readdata_from_sa;
  input   [ 31: 0] performance_counter_0_control_slave_readdata_from_sa;
  input            reset_n;
  input   [ 15: 0] sram_0_avalon_sram_slave_readdata_from_sa;
  input   [ 31: 0] sysid_control_slave_readdata_from_sa;
  input   [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] cpu_2_data_master_address_last_time;
  wire    [ 24: 0] cpu_2_data_master_address_to_slave;
  reg     [  3: 0] cpu_2_data_master_byteenable_last_time;
  reg     [  1: 0] cpu_2_data_master_dbs_address;
  wire    [  1: 0] cpu_2_data_master_dbs_increment;
  reg     [  1: 0] cpu_2_data_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_2_data_master_dbs_rdv_counter_inc;
  wire    [ 15: 0] cpu_2_data_master_dbs_write_16;
  wire    [  7: 0] cpu_2_data_master_dbs_write_8;
  wire    [ 31: 0] cpu_2_data_master_irq;
  wire             cpu_2_data_master_is_granted_some_slave;
  reg              cpu_2_data_master_latency_counter;
  wire    [  1: 0] cpu_2_data_master_next_dbs_rdv_counter;
  reg              cpu_2_data_master_read_but_no_slave_selected;
  reg              cpu_2_data_master_read_last_time;
  wire    [ 31: 0] cpu_2_data_master_readdata;
  wire             cpu_2_data_master_readdatavalid;
  wire             cpu_2_data_master_run;
  wire             cpu_2_data_master_waitrequest;
  reg              cpu_2_data_master_write_last_time;
  reg     [ 31: 0] cpu_2_data_master_writedata_last_time;
  reg     [ 15: 0] dbs_16_reg_segment_0;
  reg     [  7: 0] dbs_8_reg_segment_0;
  reg     [  7: 0] dbs_8_reg_segment_1;
  reg     [  7: 0] dbs_8_reg_segment_2;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire             p1_cpu_2_data_master_latency_counter;
  wire    [ 15: 0] p1_dbs_16_reg_segment_0;
  wire    [  7: 0] p1_dbs_8_reg_segment_0;
  wire    [  7: 0] p1_dbs_8_reg_segment_1;
  wire    [  7: 0] p1_dbs_8_reg_segment_2;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_2_data_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  wire             r_3;
  wire             r_4;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module | ~cpu_2_data_master_requests_cpu_2_jtag_debug_module) & (cpu_2_data_master_granted_cpu_2_jtag_debug_module | ~cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module) & ((~cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module | ~cpu_2_data_master_read | (1 & ~d1_cpu_2_jtag_debug_module_end_xfer & cpu_2_data_master_read))) & ((~cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module | ~cpu_2_data_master_write | (1 & cpu_2_data_master_write))) & 1 & (cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave | ~cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave) & ((~cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & ~jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa & (cpu_2_data_master_read | cpu_2_data_master_write)))) & ((~cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & ~jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa & (cpu_2_data_master_read | cpu_2_data_master_write)))) & 1 & (cpu_2_data_master_qualified_request_keys_s1 | ~cpu_2_data_master_requests_keys_s1) & (cpu_2_data_master_granted_keys_s1 | ~cpu_2_data_master_qualified_request_keys_s1) & ((~cpu_2_data_master_qualified_request_keys_s1 | ~cpu_2_data_master_read | (1 & ~d1_keys_s1_end_xfer & cpu_2_data_master_read))) & ((~cpu_2_data_master_qualified_request_keys_s1 | ~cpu_2_data_master_write | (1 & cpu_2_data_master_write))) & 1 & (cpu_2_data_master_qualified_request_mailbox_0_s1 | ~cpu_2_data_master_requests_mailbox_0_s1) & (cpu_2_data_master_granted_mailbox_0_s1 | ~cpu_2_data_master_qualified_request_mailbox_0_s1) & ((~cpu_2_data_master_qualified_request_mailbox_0_s1 | ~cpu_2_data_master_read | (1 & ~d1_mailbox_0_s1_end_xfer & cpu_2_data_master_read))) & ((~cpu_2_data_master_qualified_request_mailbox_0_s1 | ~cpu_2_data_master_write | (1 & cpu_2_data_master_write)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_2_data_master_run = r_0 & r_1 & r_2 & r_3 & r_4;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_2_data_master_qualified_request_mailbox_1_s1 | ~cpu_2_data_master_requests_mailbox_1_s1) & (cpu_2_data_master_granted_mailbox_1_s1 | ~cpu_2_data_master_qualified_request_mailbox_1_s1) & ((~cpu_2_data_master_qualified_request_mailbox_1_s1 | ~cpu_2_data_master_read | (1 & ~d1_mailbox_1_s1_end_xfer & cpu_2_data_master_read))) & ((~cpu_2_data_master_qualified_request_mailbox_1_s1 | ~cpu_2_data_master_write | (1 & cpu_2_data_master_write))) & 1 & (cpu_2_data_master_qualified_request_mailbox_2_s1 | ~cpu_2_data_master_requests_mailbox_2_s1) & (cpu_2_data_master_granted_mailbox_2_s1 | ~cpu_2_data_master_qualified_request_mailbox_2_s1) & ((~cpu_2_data_master_qualified_request_mailbox_2_s1 | ~cpu_2_data_master_read | (1 & ~d1_mailbox_2_s1_end_xfer & cpu_2_data_master_read))) & ((~cpu_2_data_master_qualified_request_mailbox_2_s1 | ~cpu_2_data_master_write | (1 & cpu_2_data_master_write))) & 1 & (cpu_2_data_master_qualified_request_mailbox_3_s1 | ~cpu_2_data_master_requests_mailbox_3_s1) & (cpu_2_data_master_granted_mailbox_3_s1 | ~cpu_2_data_master_qualified_request_mailbox_3_s1) & ((~cpu_2_data_master_qualified_request_mailbox_3_s1 | ~cpu_2_data_master_read | (1 & ~d1_mailbox_3_s1_end_xfer & cpu_2_data_master_read))) & ((~cpu_2_data_master_qualified_request_mailbox_3_s1 | ~cpu_2_data_master_write | (1 & cpu_2_data_master_write))) & 1 & ((cpu_2_data_master_qualified_request_nios_system_clock_10_in | ((cpu_2_data_master_write & !cpu_2_data_master_byteenable_nios_system_clock_10_in & cpu_2_data_master_dbs_address[1] & cpu_2_data_master_dbs_address[0])) | ~cpu_2_data_master_requests_nios_system_clock_10_in)) & ((~cpu_2_data_master_qualified_request_nios_system_clock_10_in | ~cpu_2_data_master_read | (1 & ~nios_system_clock_10_in_waitrequest_from_sa & (cpu_2_data_master_dbs_address[1] & cpu_2_data_master_dbs_address[0]) & cpu_2_data_master_read))) & ((~cpu_2_data_master_qualified_request_nios_system_clock_10_in | ~cpu_2_data_master_write | (1 & ~nios_system_clock_10_in_waitrequest_from_sa & (cpu_2_data_master_dbs_address[1] & cpu_2_data_master_dbs_address[0]) & cpu_2_data_master_write))) & 1;

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = (cpu_2_data_master_qualified_request_nios_system_clock_5_in | (cpu_2_data_master_write & !cpu_2_data_master_byteenable_nios_system_clock_5_in & cpu_2_data_master_dbs_address[1]) | ~cpu_2_data_master_requests_nios_system_clock_5_in) & ((~cpu_2_data_master_qualified_request_nios_system_clock_5_in | ~cpu_2_data_master_read | (1 & ~nios_system_clock_5_in_waitrequest_from_sa & (cpu_2_data_master_dbs_address[1]) & cpu_2_data_master_read))) & ((~cpu_2_data_master_qualified_request_nios_system_clock_5_in | ~cpu_2_data_master_write | (1 & ~nios_system_clock_5_in_waitrequest_from_sa & (cpu_2_data_master_dbs_address[1]) & cpu_2_data_master_write))) & 1 & (cpu_2_data_master_qualified_request_onchip_memory2_0_s1 | ~cpu_2_data_master_requests_onchip_memory2_0_s1) & (cpu_2_data_master_granted_onchip_memory2_0_s1 | ~cpu_2_data_master_qualified_request_onchip_memory2_0_s1) & ((~cpu_2_data_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write)))) & ((~cpu_2_data_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write)))) & 1 & (cpu_2_data_master_qualified_request_onchip_memory2_1_s1 | ~cpu_2_data_master_requests_onchip_memory2_1_s1) & (cpu_2_data_master_granted_onchip_memory2_1_s1 | ~cpu_2_data_master_qualified_request_onchip_memory2_1_s1) & ((~cpu_2_data_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write)))) & ((~cpu_2_data_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write)))) & 1 & (cpu_2_data_master_qualified_request_onchip_memory2_2_s1 | ~cpu_2_data_master_requests_onchip_memory2_2_s1) & (cpu_2_data_master_granted_onchip_memory2_2_s1 | ~cpu_2_data_master_qualified_request_onchip_memory2_2_s1) & ((~cpu_2_data_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write)))) & ((~cpu_2_data_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write))));

  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (cpu_2_data_master_qualified_request_onchip_memory2_3_s1 | ~cpu_2_data_master_requests_onchip_memory2_3_s1) & (cpu_2_data_master_granted_onchip_memory2_3_s1 | ~cpu_2_data_master_qualified_request_onchip_memory2_3_s1) & ((~cpu_2_data_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write)))) & ((~cpu_2_data_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write)))) & 1 & (cpu_2_data_master_qualified_request_performance_counter_0_control_slave | ~cpu_2_data_master_requests_performance_counter_0_control_slave) & (cpu_2_data_master_granted_performance_counter_0_control_slave | ~cpu_2_data_master_qualified_request_performance_counter_0_control_slave) & ((~cpu_2_data_master_qualified_request_performance_counter_0_control_slave | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write)))) & ((~cpu_2_data_master_qualified_request_performance_counter_0_control_slave | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write)))) & 1 & (cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave | (cpu_2_data_master_write & !cpu_2_data_master_byteenable_sram_0_avalon_sram_slave & cpu_2_data_master_dbs_address[1]) | ~cpu_2_data_master_requests_sram_0_avalon_sram_slave) & (cpu_2_data_master_granted_sram_0_avalon_sram_slave | ~cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave) & ((~cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_2_data_master_read | (1 & (cpu_2_data_master_dbs_address[1]) & cpu_2_data_master_read))) & ((~cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_2_data_master_write | (1 & (cpu_2_data_master_dbs_address[1]) & cpu_2_data_master_write))) & 1 & (cpu_2_data_master_qualified_request_sysid_control_slave | ~cpu_2_data_master_requests_sysid_control_slave) & (cpu_2_data_master_granted_sysid_control_slave | ~cpu_2_data_master_qualified_request_sysid_control_slave) & ((~cpu_2_data_master_qualified_request_sysid_control_slave | ~cpu_2_data_master_read | (1 & ~d1_sysid_control_slave_end_xfer & cpu_2_data_master_read)));

  //r_4 master_run cascaded wait assignment, which is an e_assign
  assign r_4 = ((~cpu_2_data_master_qualified_request_sysid_control_slave | ~cpu_2_data_master_write | (1 & cpu_2_data_master_write))) & 1 & (cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) & (cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave | ~cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave) & ((~cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write)))) & ((~cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~(cpu_2_data_master_read | cpu_2_data_master_write) | (1 & (cpu_2_data_master_read | cpu_2_data_master_write))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_2_data_master_address_to_slave = cpu_2_data_master_address[24 : 0];

  //cpu_2_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_read_but_no_slave_selected <= 0;
      else 
        cpu_2_data_master_read_but_no_slave_selected <= cpu_2_data_master_read & cpu_2_data_master_run & ~cpu_2_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_2_data_master_is_granted_some_slave = cpu_2_data_master_granted_cpu_2_jtag_debug_module |
    cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave |
    cpu_2_data_master_granted_keys_s1 |
    cpu_2_data_master_granted_mailbox_0_s1 |
    cpu_2_data_master_granted_mailbox_1_s1 |
    cpu_2_data_master_granted_mailbox_2_s1 |
    cpu_2_data_master_granted_mailbox_3_s1 |
    cpu_2_data_master_granted_nios_system_clock_10_in |
    cpu_2_data_master_granted_nios_system_clock_5_in |
    cpu_2_data_master_granted_onchip_memory2_0_s1 |
    cpu_2_data_master_granted_onchip_memory2_1_s1 |
    cpu_2_data_master_granted_onchip_memory2_2_s1 |
    cpu_2_data_master_granted_onchip_memory2_3_s1 |
    cpu_2_data_master_granted_performance_counter_0_control_slave |
    cpu_2_data_master_granted_sram_0_avalon_sram_slave |
    cpu_2_data_master_granted_sysid_control_slave |
    cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_2_data_master_readdatavalid = cpu_2_data_master_read_data_valid_onchip_memory2_0_s1 |
    cpu_2_data_master_read_data_valid_onchip_memory2_1_s1 |
    cpu_2_data_master_read_data_valid_onchip_memory2_2_s1 |
    cpu_2_data_master_read_data_valid_onchip_memory2_3_s1 |
    cpu_2_data_master_read_data_valid_performance_counter_0_control_slave |
    (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave & dbs_rdv_counter_overflow) |
    cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_2_data_master_readdatavalid = cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_data_valid_keys_s1 |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_data_valid_mailbox_0_s1 |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_data_valid_mailbox_1_s1 |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_data_valid_mailbox_2_s1 |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_data_valid_mailbox_3_s1 |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    (cpu_2_data_master_read_data_valid_nios_system_clock_10_in & dbs_counter_overflow) |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    (cpu_2_data_master_read_data_valid_nios_system_clock_5_in & dbs_counter_overflow) |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid |
    cpu_2_data_master_read_data_valid_sysid_control_slave |
    cpu_2_data_master_read_but_no_slave_selected |
    pre_flush_cpu_2_data_master_readdatavalid;

  //cpu_2/data_master readdata mux, which is an e_mux
  assign cpu_2_data_master_readdata = ({32 {~(cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module & cpu_2_data_master_read)}} | cpu_2_jtag_debug_module_readdata_from_sa) &
    ({32 {~(cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave & cpu_2_data_master_read)}} | jtag_uart_2_avalon_jtag_slave_readdata_from_sa) &
    ({32 {~(cpu_2_data_master_qualified_request_keys_s1 & cpu_2_data_master_read)}} | keys_s1_readdata_from_sa) &
    ({32 {~(cpu_2_data_master_qualified_request_mailbox_0_s1 & cpu_2_data_master_read)}} | mailbox_0_s1_readdata_from_sa) &
    ({32 {~(cpu_2_data_master_qualified_request_mailbox_1_s1 & cpu_2_data_master_read)}} | mailbox_1_s1_readdata_from_sa) &
    ({32 {~(cpu_2_data_master_qualified_request_mailbox_2_s1 & cpu_2_data_master_read)}} | mailbox_2_s1_readdata_from_sa) &
    ({32 {~(cpu_2_data_master_qualified_request_mailbox_3_s1 & cpu_2_data_master_read)}} | mailbox_3_s1_readdata_from_sa) &
    ({32 {~(cpu_2_data_master_qualified_request_nios_system_clock_10_in & cpu_2_data_master_read)}} | {nios_system_clock_10_in_readdata_from_sa[7 : 0],
    dbs_8_reg_segment_2,
    dbs_8_reg_segment_1,
    dbs_8_reg_segment_0}) &
    ({32 {~(cpu_2_data_master_qualified_request_nios_system_clock_5_in & cpu_2_data_master_read)}} | {nios_system_clock_5_in_readdata_from_sa[15 : 0],
    dbs_16_reg_segment_0}) &
    ({32 {~cpu_2_data_master_read_data_valid_onchip_memory2_0_s1}} | onchip_memory2_0_s1_readdata_from_sa) &
    ({32 {~cpu_2_data_master_read_data_valid_onchip_memory2_1_s1}} | onchip_memory2_1_s1_readdata_from_sa) &
    ({32 {~cpu_2_data_master_read_data_valid_onchip_memory2_2_s1}} | onchip_memory2_2_s1_readdata_from_sa) &
    ({32 {~cpu_2_data_master_read_data_valid_onchip_memory2_3_s1}} | onchip_memory2_3_s1_readdata_from_sa) &
    ({32 {~cpu_2_data_master_read_data_valid_performance_counter_0_control_slave}} | performance_counter_0_control_slave_readdata_from_sa) &
    ({32 {~cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave}} | {sram_0_avalon_sram_slave_readdata_from_sa[15 : 0],
    dbs_latent_16_reg_segment_0}) &
    ({32 {~(cpu_2_data_master_qualified_request_sysid_control_slave & cpu_2_data_master_read)}} | sysid_control_slave_readdata_from_sa) &
    ({32 {~cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave}} | video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_2_data_master_waitrequest = ~cpu_2_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_latency_counter <= 0;
      else 
        cpu_2_data_master_latency_counter <= p1_cpu_2_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_2_data_master_latency_counter = ((cpu_2_data_master_run & cpu_2_data_master_read))? latency_load_value :
    (cpu_2_data_master_latency_counter)? cpu_2_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({1 {cpu_2_data_master_requests_onchip_memory2_0_s1}} & 1) |
    ({1 {cpu_2_data_master_requests_onchip_memory2_1_s1}} & 1) |
    ({1 {cpu_2_data_master_requests_onchip_memory2_2_s1}} & 1) |
    ({1 {cpu_2_data_master_requests_onchip_memory2_3_s1}} & 1) |
    ({1 {cpu_2_data_master_requests_performance_counter_0_control_slave}} & 1) |
    ({1 {cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave}} & 1);

  //irq assign, which is an e_assign
  assign cpu_2_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    jtag_uart_2_avalon_jtag_slave_irq_from_sa,
    1'b0};

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (((~0) & cpu_2_data_master_requests_nios_system_clock_10_in & cpu_2_data_master_write & !cpu_2_data_master_byteenable_nios_system_clock_10_in)) |
    (cpu_2_data_master_granted_nios_system_clock_10_in & cpu_2_data_master_read & 1 & 1 & ~nios_system_clock_10_in_waitrequest_from_sa) |
    (cpu_2_data_master_granted_nios_system_clock_10_in & cpu_2_data_master_write & 1 & 1 & ~nios_system_clock_10_in_waitrequest_from_sa) |
    (((~0) & cpu_2_data_master_requests_nios_system_clock_5_in & cpu_2_data_master_write & !cpu_2_data_master_byteenable_nios_system_clock_5_in)) |
    (cpu_2_data_master_granted_nios_system_clock_5_in & cpu_2_data_master_read & 1 & 1 & ~nios_system_clock_5_in_waitrequest_from_sa) |
    (cpu_2_data_master_granted_nios_system_clock_5_in & cpu_2_data_master_write & 1 & 1 & ~nios_system_clock_5_in_waitrequest_from_sa) |
    (((~0) & cpu_2_data_master_requests_sram_0_avalon_sram_slave & cpu_2_data_master_write & !cpu_2_data_master_byteenable_sram_0_avalon_sram_slave)) |
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave & cpu_2_data_master_read & 1 & 1) |
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave & cpu_2_data_master_write & 1 & 1);

  //input to dbs-8 stored 0, which is an e_mux
  assign p1_dbs_8_reg_segment_0 = nios_system_clock_10_in_readdata_from_sa;

  //dbs register for dbs-8 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_2_data_master_dbs_address[1 : 0]) == 0))
          dbs_8_reg_segment_0 <= p1_dbs_8_reg_segment_0;
    end


  //input to dbs-8 stored 1, which is an e_mux
  assign p1_dbs_8_reg_segment_1 = nios_system_clock_10_in_readdata_from_sa;

  //dbs register for dbs-8 segment 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_1 <= 0;
      else if (dbs_count_enable & ((cpu_2_data_master_dbs_address[1 : 0]) == 1))
          dbs_8_reg_segment_1 <= p1_dbs_8_reg_segment_1;
    end


  //input to dbs-8 stored 2, which is an e_mux
  assign p1_dbs_8_reg_segment_2 = nios_system_clock_10_in_readdata_from_sa;

  //dbs register for dbs-8 segment 2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_2 <= 0;
      else if (dbs_count_enable & ((cpu_2_data_master_dbs_address[1 : 0]) == 2))
          dbs_8_reg_segment_2 <= p1_dbs_8_reg_segment_2;
    end


  //mux write dbs 2, which is an e_mux
  assign cpu_2_data_master_dbs_write_8 = ((cpu_2_data_master_dbs_address[1 : 0] == 0))? cpu_2_data_master_writedata[7 : 0] :
    ((cpu_2_data_master_dbs_address[1 : 0] == 1))? cpu_2_data_master_writedata[15 : 8] :
    ((cpu_2_data_master_dbs_address[1 : 0] == 2))? cpu_2_data_master_writedata[23 : 16] :
    cpu_2_data_master_writedata[31 : 24];

  //dbs count increment, which is an e_mux
  assign cpu_2_data_master_dbs_increment = (cpu_2_data_master_requests_nios_system_clock_10_in)? 1 :
    (cpu_2_data_master_requests_nios_system_clock_5_in)? 2 :
    (cpu_2_data_master_requests_sram_0_avalon_sram_slave)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_2_data_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_2_data_master_dbs_address + cpu_2_data_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_2_data_master_dbs_address <= next_dbs_address;
    end


  //input to dbs-16 stored 0, which is an e_mux
  assign p1_dbs_16_reg_segment_0 = nios_system_clock_5_in_readdata_from_sa;

  //dbs register for dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_16_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_2_data_master_dbs_address[1]) == 0))
          dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
    end


  //mux write dbs 1, which is an e_mux
  assign cpu_2_data_master_dbs_write_16 = (cpu_2_data_master_dbs_address[1])? cpu_2_data_master_writedata[31 : 16] :
    (~(cpu_2_data_master_dbs_address[1]))? cpu_2_data_master_writedata[15 : 0] :
    (cpu_2_data_master_dbs_address[1])? cpu_2_data_master_writedata[31 : 16] :
    cpu_2_data_master_writedata[15 : 0];

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = sram_0_avalon_sram_slave_readdata_from_sa;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_2_data_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_2_data_master_next_dbs_rdv_counter = cpu_2_data_master_dbs_rdv_counter + cpu_2_data_master_dbs_rdv_counter_inc;

  //cpu_2_data_master_rdv_inc_mux, which is an e_mux
  assign cpu_2_data_master_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_2_data_master_dbs_rdv_counter <= cpu_2_data_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_2_data_master_dbs_rdv_counter[1] & ~cpu_2_data_master_next_dbs_rdv_counter[1];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_2_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_address_last_time <= 0;
      else 
        cpu_2_data_master_address_last_time <= cpu_2_data_master_address;
    end


  //cpu_2/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_2_data_master_waitrequest & (cpu_2_data_master_read | cpu_2_data_master_write);
    end


  //cpu_2_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_2_data_master_address != cpu_2_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_2_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_2_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_byteenable_last_time <= 0;
      else 
        cpu_2_data_master_byteenable_last_time <= cpu_2_data_master_byteenable;
    end


  //cpu_2_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_2_data_master_byteenable != cpu_2_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_2_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_2_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_read_last_time <= 0;
      else 
        cpu_2_data_master_read_last_time <= cpu_2_data_master_read;
    end


  //cpu_2_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_2_data_master_read != cpu_2_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_2_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_2_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_write_last_time <= 0;
      else 
        cpu_2_data_master_write_last_time <= cpu_2_data_master_write;
    end


  //cpu_2_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_2_data_master_write != cpu_2_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_2_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_2_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_writedata_last_time <= 0;
      else 
        cpu_2_data_master_writedata_last_time <= cpu_2_data_master_writedata;
    end


  //cpu_2_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_2_data_master_writedata != cpu_2_data_master_writedata_last_time) & cpu_2_data_master_write)
        begin
          $write("%0d ns: cpu_2_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_2_instruction_master_arbitrator (
                                             // inputs:
                                              clk,
                                              cpu_2_instruction_master_address,
                                              cpu_2_instruction_master_granted_cpu_2_jtag_debug_module,
                                              cpu_2_instruction_master_granted_nios_system_clock_4_in,
                                              cpu_2_instruction_master_granted_onchip_memory2_0_s1,
                                              cpu_2_instruction_master_granted_onchip_memory2_1_s1,
                                              cpu_2_instruction_master_granted_onchip_memory2_2_s1,
                                              cpu_2_instruction_master_granted_onchip_memory2_3_s1,
                                              cpu_2_instruction_master_granted_sram_0_avalon_sram_slave,
                                              cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module,
                                              cpu_2_instruction_master_qualified_request_nios_system_clock_4_in,
                                              cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1,
                                              cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1,
                                              cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1,
                                              cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1,
                                              cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave,
                                              cpu_2_instruction_master_read,
                                              cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module,
                                              cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in,
                                              cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1,
                                              cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1,
                                              cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1,
                                              cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1,
                                              cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave,
                                              cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                              cpu_2_instruction_master_requests_cpu_2_jtag_debug_module,
                                              cpu_2_instruction_master_requests_nios_system_clock_4_in,
                                              cpu_2_instruction_master_requests_onchip_memory2_0_s1,
                                              cpu_2_instruction_master_requests_onchip_memory2_1_s1,
                                              cpu_2_instruction_master_requests_onchip_memory2_2_s1,
                                              cpu_2_instruction_master_requests_onchip_memory2_3_s1,
                                              cpu_2_instruction_master_requests_sram_0_avalon_sram_slave,
                                              cpu_2_jtag_debug_module_readdata_from_sa,
                                              d1_cpu_2_jtag_debug_module_end_xfer,
                                              d1_nios_system_clock_4_in_end_xfer,
                                              d1_onchip_memory2_0_s1_end_xfer,
                                              d1_onchip_memory2_1_s1_end_xfer,
                                              d1_onchip_memory2_2_s1_end_xfer,
                                              d1_onchip_memory2_3_s1_end_xfer,
                                              d1_sram_0_avalon_sram_slave_end_xfer,
                                              nios_system_clock_4_in_readdata_from_sa,
                                              nios_system_clock_4_in_waitrequest_from_sa,
                                              onchip_memory2_0_s1_readdata_from_sa,
                                              onchip_memory2_1_s1_readdata_from_sa,
                                              onchip_memory2_2_s1_readdata_from_sa,
                                              onchip_memory2_3_s1_readdata_from_sa,
                                              reset_n,
                                              sram_0_avalon_sram_slave_readdata_from_sa,

                                             // outputs:
                                              cpu_2_instruction_master_address_to_slave,
                                              cpu_2_instruction_master_dbs_address,
                                              cpu_2_instruction_master_latency_counter,
                                              cpu_2_instruction_master_readdata,
                                              cpu_2_instruction_master_readdatavalid,
                                              cpu_2_instruction_master_waitrequest
                                           )
;

  output  [ 24: 0] cpu_2_instruction_master_address_to_slave;
  output  [  1: 0] cpu_2_instruction_master_dbs_address;
  output           cpu_2_instruction_master_latency_counter;
  output  [ 31: 0] cpu_2_instruction_master_readdata;
  output           cpu_2_instruction_master_readdatavalid;
  output           cpu_2_instruction_master_waitrequest;
  input            clk;
  input   [ 24: 0] cpu_2_instruction_master_address;
  input            cpu_2_instruction_master_granted_cpu_2_jtag_debug_module;
  input            cpu_2_instruction_master_granted_nios_system_clock_4_in;
  input            cpu_2_instruction_master_granted_onchip_memory2_0_s1;
  input            cpu_2_instruction_master_granted_onchip_memory2_1_s1;
  input            cpu_2_instruction_master_granted_onchip_memory2_2_s1;
  input            cpu_2_instruction_master_granted_onchip_memory2_3_s1;
  input            cpu_2_instruction_master_granted_sram_0_avalon_sram_slave;
  input            cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module;
  input            cpu_2_instruction_master_qualified_request_nios_system_clock_4_in;
  input            cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1;
  input            cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1;
  input            cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1;
  input            cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1;
  input            cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  input            cpu_2_instruction_master_read;
  input            cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module;
  input            cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in;
  input            cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1;
  input            cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1;
  input            cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1;
  input            cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1;
  input            cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  input            cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_instruction_master_requests_cpu_2_jtag_debug_module;
  input            cpu_2_instruction_master_requests_nios_system_clock_4_in;
  input            cpu_2_instruction_master_requests_onchip_memory2_0_s1;
  input            cpu_2_instruction_master_requests_onchip_memory2_1_s1;
  input            cpu_2_instruction_master_requests_onchip_memory2_2_s1;
  input            cpu_2_instruction_master_requests_onchip_memory2_3_s1;
  input            cpu_2_instruction_master_requests_sram_0_avalon_sram_slave;
  input   [ 31: 0] cpu_2_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_2_jtag_debug_module_end_xfer;
  input            d1_nios_system_clock_4_in_end_xfer;
  input            d1_onchip_memory2_0_s1_end_xfer;
  input            d1_onchip_memory2_1_s1_end_xfer;
  input            d1_onchip_memory2_2_s1_end_xfer;
  input            d1_onchip_memory2_3_s1_end_xfer;
  input            d1_sram_0_avalon_sram_slave_end_xfer;
  input   [ 15: 0] nios_system_clock_4_in_readdata_from_sa;
  input            nios_system_clock_4_in_waitrequest_from_sa;
  input   [ 31: 0] onchip_memory2_0_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_1_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_2_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_3_s1_readdata_from_sa;
  input            reset_n;
  input   [ 15: 0] sram_0_avalon_sram_slave_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] cpu_2_instruction_master_address_last_time;
  wire    [ 24: 0] cpu_2_instruction_master_address_to_slave;
  reg     [  1: 0] cpu_2_instruction_master_dbs_address;
  wire    [  1: 0] cpu_2_instruction_master_dbs_increment;
  reg     [  1: 0] cpu_2_instruction_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_2_instruction_master_dbs_rdv_counter_inc;
  wire             cpu_2_instruction_master_is_granted_some_slave;
  reg              cpu_2_instruction_master_latency_counter;
  wire    [  1: 0] cpu_2_instruction_master_next_dbs_rdv_counter;
  reg              cpu_2_instruction_master_read_but_no_slave_selected;
  reg              cpu_2_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_2_instruction_master_readdata;
  wire             cpu_2_instruction_master_readdatavalid;
  wire             cpu_2_instruction_master_run;
  wire             cpu_2_instruction_master_waitrequest;
  reg     [ 15: 0] dbs_16_reg_segment_0;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire             p1_cpu_2_instruction_master_latency_counter;
  wire    [ 15: 0] p1_dbs_16_reg_segment_0;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_2_instruction_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  wire             r_3;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module | ~cpu_2_instruction_master_requests_cpu_2_jtag_debug_module) & (cpu_2_instruction_master_granted_cpu_2_jtag_debug_module | ~cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module) & ((~cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module | ~cpu_2_instruction_master_read | (1 & ~d1_cpu_2_jtag_debug_module_end_xfer & cpu_2_instruction_master_read)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_2_instruction_master_run = r_0 & r_1 & r_2 & r_3;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_2_instruction_master_qualified_request_nios_system_clock_4_in | ~cpu_2_instruction_master_requests_nios_system_clock_4_in) & ((~cpu_2_instruction_master_qualified_request_nios_system_clock_4_in | ~cpu_2_instruction_master_read | (1 & ~nios_system_clock_4_in_waitrequest_from_sa & (cpu_2_instruction_master_dbs_address[1]) & cpu_2_instruction_master_read)));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1 | ~cpu_2_instruction_master_requests_onchip_memory2_0_s1) & (cpu_2_instruction_master_granted_onchip_memory2_0_s1 | ~cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1) & ((~cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_2_instruction_master_read) | (1 & (cpu_2_instruction_master_read)))) & 1 & (cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1 | ~cpu_2_instruction_master_requests_onchip_memory2_1_s1) & (cpu_2_instruction_master_granted_onchip_memory2_1_s1 | ~cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1) & ((~cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_2_instruction_master_read) | (1 & (cpu_2_instruction_master_read)))) & 1 & (cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1 | ~cpu_2_instruction_master_requests_onchip_memory2_2_s1) & (cpu_2_instruction_master_granted_onchip_memory2_2_s1 | ~cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1) & ((~cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_2_instruction_master_read) | (1 & (cpu_2_instruction_master_read))));

  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1 | ~cpu_2_instruction_master_requests_onchip_memory2_3_s1) & (cpu_2_instruction_master_granted_onchip_memory2_3_s1 | ~cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1) & ((~cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_2_instruction_master_read) | (1 & (cpu_2_instruction_master_read)))) & 1 & (cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_2_instruction_master_requests_sram_0_avalon_sram_slave) & (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave | ~cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave) & ((~cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_2_instruction_master_read | (1 & (cpu_2_instruction_master_dbs_address[1]) & cpu_2_instruction_master_read)));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_2_instruction_master_address_to_slave = cpu_2_instruction_master_address[24 : 0];

  //cpu_2_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_2_instruction_master_read_but_no_slave_selected <= cpu_2_instruction_master_read & cpu_2_instruction_master_run & ~cpu_2_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_2_instruction_master_is_granted_some_slave = cpu_2_instruction_master_granted_cpu_2_jtag_debug_module |
    cpu_2_instruction_master_granted_nios_system_clock_4_in |
    cpu_2_instruction_master_granted_onchip_memory2_0_s1 |
    cpu_2_instruction_master_granted_onchip_memory2_1_s1 |
    cpu_2_instruction_master_granted_onchip_memory2_2_s1 |
    cpu_2_instruction_master_granted_onchip_memory2_3_s1 |
    cpu_2_instruction_master_granted_sram_0_avalon_sram_slave;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_2_instruction_master_readdatavalid = cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1 |
    cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1 |
    cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1 |
    cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1 |
    (cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave & dbs_rdv_counter_overflow);

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_2_instruction_master_readdatavalid = cpu_2_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_2_instruction_master_readdatavalid |
    cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module |
    cpu_2_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_2_instruction_master_readdatavalid |
    (cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in & dbs_counter_overflow) |
    cpu_2_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_2_instruction_master_readdatavalid |
    cpu_2_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_2_instruction_master_readdatavalid |
    cpu_2_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_2_instruction_master_readdatavalid |
    cpu_2_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_2_instruction_master_readdatavalid |
    cpu_2_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_2_instruction_master_readdatavalid;

  //cpu_2/instruction_master readdata mux, which is an e_mux
  assign cpu_2_instruction_master_readdata = ({32 {~(cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module & cpu_2_instruction_master_read)}} | cpu_2_jtag_debug_module_readdata_from_sa) &
    ({32 {~(cpu_2_instruction_master_qualified_request_nios_system_clock_4_in & cpu_2_instruction_master_read)}} | {nios_system_clock_4_in_readdata_from_sa[15 : 0],
    dbs_16_reg_segment_0}) &
    ({32 {~cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1}} | onchip_memory2_0_s1_readdata_from_sa) &
    ({32 {~cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1}} | onchip_memory2_1_s1_readdata_from_sa) &
    ({32 {~cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1}} | onchip_memory2_2_s1_readdata_from_sa) &
    ({32 {~cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1}} | onchip_memory2_3_s1_readdata_from_sa) &
    ({32 {~cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave}} | {sram_0_avalon_sram_slave_readdata_from_sa[15 : 0],
    dbs_latent_16_reg_segment_0});

  //actual waitrequest port, which is an e_assign
  assign cpu_2_instruction_master_waitrequest = ~cpu_2_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_instruction_master_latency_counter <= 0;
      else 
        cpu_2_instruction_master_latency_counter <= p1_cpu_2_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_2_instruction_master_latency_counter = ((cpu_2_instruction_master_run & cpu_2_instruction_master_read))? latency_load_value :
    (cpu_2_instruction_master_latency_counter)? cpu_2_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({1 {cpu_2_instruction_master_requests_onchip_memory2_0_s1}} & 1) |
    ({1 {cpu_2_instruction_master_requests_onchip_memory2_1_s1}} & 1) |
    ({1 {cpu_2_instruction_master_requests_onchip_memory2_2_s1}} & 1) |
    ({1 {cpu_2_instruction_master_requests_onchip_memory2_3_s1}} & 1);

  //input to dbs-16 stored 0, which is an e_mux
  assign p1_dbs_16_reg_segment_0 = nios_system_clock_4_in_readdata_from_sa;

  //dbs register for dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_16_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_2_instruction_master_dbs_address[1]) == 0))
          dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
    end


  //dbs count increment, which is an e_mux
  assign cpu_2_instruction_master_dbs_increment = (cpu_2_instruction_master_requests_nios_system_clock_4_in)? 2 :
    (cpu_2_instruction_master_requests_sram_0_avalon_sram_slave)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_2_instruction_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_2_instruction_master_dbs_address + cpu_2_instruction_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_instruction_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_2_instruction_master_dbs_address <= next_dbs_address;
    end


  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (cpu_2_instruction_master_granted_nios_system_clock_4_in & cpu_2_instruction_master_read & 1 & 1 & ~nios_system_clock_4_in_waitrequest_from_sa) |
    (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave & cpu_2_instruction_master_read & 1 & 1);

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = sram_0_avalon_sram_slave_readdata_from_sa;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_2_instruction_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_2_instruction_master_next_dbs_rdv_counter = cpu_2_instruction_master_dbs_rdv_counter + cpu_2_instruction_master_dbs_rdv_counter_inc;

  //cpu_2_instruction_master_rdv_inc_mux, which is an e_mux
  assign cpu_2_instruction_master_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_instruction_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_2_instruction_master_dbs_rdv_counter <= cpu_2_instruction_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_2_instruction_master_dbs_rdv_counter[1] & ~cpu_2_instruction_master_next_dbs_rdv_counter[1];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_2_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_instruction_master_address_last_time <= 0;
      else 
        cpu_2_instruction_master_address_last_time <= cpu_2_instruction_master_address;
    end


  //cpu_2/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_2_instruction_master_waitrequest & (cpu_2_instruction_master_read);
    end


  //cpu_2_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_2_instruction_master_address != cpu_2_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_2_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_2_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_instruction_master_read_last_time <= 0;
      else 
        cpu_2_instruction_master_read_last_time <= cpu_2_instruction_master_read;
    end


  //cpu_2_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_2_instruction_master_read != cpu_2_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_2_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_2_altera_nios_custom_instr_floating_point_inst_s1_arbitrator (
                                                                          // inputs:
                                                                           clk,
                                                                           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done,
                                                                           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result,
                                                                           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select,
                                                                           cpu_2_custom_instruction_master_multi_clk_en,
                                                                           cpu_2_custom_instruction_master_multi_dataa,
                                                                           cpu_2_custom_instruction_master_multi_datab,
                                                                           cpu_2_custom_instruction_master_multi_n,
                                                                           cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1,
                                                                           reset_n,

                                                                          // outputs:
                                                                           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_clk_en,
                                                                           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_dataa,
                                                                           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_datab,
                                                                           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa,
                                                                           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_n,
                                                                           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_reset,
                                                                           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa,
                                                                           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_start
                                                                        )
;

  output           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  output  [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  output  [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_datab;
  output           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  output  [  1: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_n;
  output           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_reset;
  output  [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  output           cpu_2_altera_nios_custom_instr_floating_point_inst_s1_start;
  input            clk;
  input            cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done;
  input   [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result;
  input            cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select;
  input            cpu_2_custom_instruction_master_multi_clk_en;
  input   [ 31: 0] cpu_2_custom_instruction_master_multi_dataa;
  input   [ 31: 0] cpu_2_custom_instruction_master_multi_datab;
  input   [  7: 0] cpu_2_custom_instruction_master_multi_n;
  input            cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1;
  input            reset_n;

  wire             cpu_2_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  wire    [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  wire    [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_datab;
  wire             cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  wire    [  1: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_n;
  wire             cpu_2_altera_nios_custom_instr_floating_point_inst_s1_reset;
  wire    [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  wire             cpu_2_altera_nios_custom_instr_floating_point_inst_s1_start;
  assign cpu_2_altera_nios_custom_instr_floating_point_inst_s1_clk_en = cpu_2_custom_instruction_master_multi_clk_en;
  assign cpu_2_altera_nios_custom_instr_floating_point_inst_s1_dataa = cpu_2_custom_instruction_master_multi_dataa;
  assign cpu_2_altera_nios_custom_instr_floating_point_inst_s1_datab = cpu_2_custom_instruction_master_multi_datab;
  assign cpu_2_altera_nios_custom_instr_floating_point_inst_s1_n = cpu_2_custom_instruction_master_multi_n;
  assign cpu_2_altera_nios_custom_instr_floating_point_inst_s1_start = cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1;
  //assign cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa = cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa = cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result;

  //assign cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa = cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa = cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done;

  //cpu_2_altera_nios_custom_instr_floating_point_inst/s1 local reset_n, which is an e_assign
  assign cpu_2_altera_nios_custom_instr_floating_point_inst_s1_reset = ~reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_3_jtag_debug_module_arbitrator (
                                            // inputs:
                                             clk,
                                             cpu_3_data_master_address_to_slave,
                                             cpu_3_data_master_byteenable,
                                             cpu_3_data_master_debugaccess,
                                             cpu_3_data_master_latency_counter,
                                             cpu_3_data_master_read,
                                             cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                             cpu_3_data_master_write,
                                             cpu_3_data_master_writedata,
                                             cpu_3_instruction_master_address_to_slave,
                                             cpu_3_instruction_master_latency_counter,
                                             cpu_3_instruction_master_read,
                                             cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                             cpu_3_jtag_debug_module_readdata,
                                             cpu_3_jtag_debug_module_resetrequest,
                                             reset_n,

                                            // outputs:
                                             cpu_3_data_master_granted_cpu_3_jtag_debug_module,
                                             cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module,
                                             cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module,
                                             cpu_3_data_master_requests_cpu_3_jtag_debug_module,
                                             cpu_3_instruction_master_granted_cpu_3_jtag_debug_module,
                                             cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module,
                                             cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module,
                                             cpu_3_instruction_master_requests_cpu_3_jtag_debug_module,
                                             cpu_3_jtag_debug_module_address,
                                             cpu_3_jtag_debug_module_begintransfer,
                                             cpu_3_jtag_debug_module_byteenable,
                                             cpu_3_jtag_debug_module_chipselect,
                                             cpu_3_jtag_debug_module_debugaccess,
                                             cpu_3_jtag_debug_module_readdata_from_sa,
                                             cpu_3_jtag_debug_module_resetrequest_from_sa,
                                             cpu_3_jtag_debug_module_write,
                                             cpu_3_jtag_debug_module_writedata,
                                             d1_cpu_3_jtag_debug_module_end_xfer
                                          )
;

  output           cpu_3_data_master_granted_cpu_3_jtag_debug_module;
  output           cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module;
  output           cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module;
  output           cpu_3_data_master_requests_cpu_3_jtag_debug_module;
  output           cpu_3_instruction_master_granted_cpu_3_jtag_debug_module;
  output           cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module;
  output           cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module;
  output           cpu_3_instruction_master_requests_cpu_3_jtag_debug_module;
  output  [  8: 0] cpu_3_jtag_debug_module_address;
  output           cpu_3_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_3_jtag_debug_module_byteenable;
  output           cpu_3_jtag_debug_module_chipselect;
  output           cpu_3_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_3_jtag_debug_module_readdata_from_sa;
  output           cpu_3_jtag_debug_module_resetrequest_from_sa;
  output           cpu_3_jtag_debug_module_write;
  output  [ 31: 0] cpu_3_jtag_debug_module_writedata;
  output           d1_cpu_3_jtag_debug_module_end_xfer;
  input            clk;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input   [  3: 0] cpu_3_data_master_byteenable;
  input            cpu_3_data_master_debugaccess;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 24: 0] cpu_3_instruction_master_address_to_slave;
  input            cpu_3_instruction_master_latency_counter;
  input            cpu_3_instruction_master_read;
  input            cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 31: 0] cpu_3_jtag_debug_module_readdata;
  input            cpu_3_jtag_debug_module_resetrequest;
  input            reset_n;

  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_cpu_3_jtag_debug_module;
  wire             cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module;
  wire             cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module;
  wire             cpu_3_data_master_requests_cpu_3_jtag_debug_module;
  wire             cpu_3_data_master_saved_grant_cpu_3_jtag_debug_module;
  wire             cpu_3_instruction_master_arbiterlock;
  wire             cpu_3_instruction_master_arbiterlock2;
  wire             cpu_3_instruction_master_continuerequest;
  wire             cpu_3_instruction_master_granted_cpu_3_jtag_debug_module;
  wire             cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module;
  wire             cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module;
  wire             cpu_3_instruction_master_requests_cpu_3_jtag_debug_module;
  wire             cpu_3_instruction_master_saved_grant_cpu_3_jtag_debug_module;
  wire    [  8: 0] cpu_3_jtag_debug_module_address;
  wire             cpu_3_jtag_debug_module_allgrants;
  wire             cpu_3_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_3_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_3_jtag_debug_module_any_continuerequest;
  reg     [  1: 0] cpu_3_jtag_debug_module_arb_addend;
  wire             cpu_3_jtag_debug_module_arb_counter_enable;
  reg     [  2: 0] cpu_3_jtag_debug_module_arb_share_counter;
  wire    [  2: 0] cpu_3_jtag_debug_module_arb_share_counter_next_value;
  wire    [  2: 0] cpu_3_jtag_debug_module_arb_share_set_values;
  wire    [  1: 0] cpu_3_jtag_debug_module_arb_winner;
  wire             cpu_3_jtag_debug_module_arbitration_holdoff_internal;
  wire             cpu_3_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_3_jtag_debug_module_begins_xfer;
  wire             cpu_3_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_3_jtag_debug_module_byteenable;
  wire             cpu_3_jtag_debug_module_chipselect;
  wire    [  3: 0] cpu_3_jtag_debug_module_chosen_master_double_vector;
  wire    [  1: 0] cpu_3_jtag_debug_module_chosen_master_rot_left;
  wire             cpu_3_jtag_debug_module_debugaccess;
  wire             cpu_3_jtag_debug_module_end_xfer;
  wire             cpu_3_jtag_debug_module_firsttransfer;
  wire    [  1: 0] cpu_3_jtag_debug_module_grant_vector;
  wire             cpu_3_jtag_debug_module_in_a_read_cycle;
  wire             cpu_3_jtag_debug_module_in_a_write_cycle;
  wire    [  1: 0] cpu_3_jtag_debug_module_master_qreq_vector;
  wire             cpu_3_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_3_jtag_debug_module_readdata_from_sa;
  reg              cpu_3_jtag_debug_module_reg_firsttransfer;
  wire             cpu_3_jtag_debug_module_resetrequest_from_sa;
  reg     [  1: 0] cpu_3_jtag_debug_module_saved_chosen_master_vector;
  reg              cpu_3_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_3_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_3_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_3_jtag_debug_module_waits_for_read;
  wire             cpu_3_jtag_debug_module_waits_for_write;
  wire             cpu_3_jtag_debug_module_write;
  wire    [ 31: 0] cpu_3_jtag_debug_module_writedata;
  reg              d1_cpu_3_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_3_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_3_data_master_granted_slave_cpu_3_jtag_debug_module;
  reg              last_cycle_cpu_3_instruction_master_granted_slave_cpu_3_jtag_debug_module;
  wire    [ 24: 0] shifted_address_to_cpu_3_jtag_debug_module_from_cpu_3_data_master;
  wire    [ 24: 0] shifted_address_to_cpu_3_jtag_debug_module_from_cpu_3_instruction_master;
  wire             wait_for_cpu_3_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_3_jtag_debug_module_end_xfer;
    end


  assign cpu_3_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module | cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module));
  //assign cpu_3_jtag_debug_module_readdata_from_sa = cpu_3_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_3_jtag_debug_module_readdata_from_sa = cpu_3_jtag_debug_module_readdata;

  assign cpu_3_data_master_requests_cpu_3_jtag_debug_module = ({cpu_3_data_master_address_to_slave[24 : 11] , 11'b0} == 25'h2000) & (cpu_3_data_master_read | cpu_3_data_master_write);
  //cpu_3_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_3_jtag_debug_module_arb_share_set_values = 1;

  //cpu_3_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_3_jtag_debug_module_non_bursting_master_requests = cpu_3_data_master_requests_cpu_3_jtag_debug_module |
    cpu_3_instruction_master_requests_cpu_3_jtag_debug_module |
    cpu_3_data_master_requests_cpu_3_jtag_debug_module |
    cpu_3_instruction_master_requests_cpu_3_jtag_debug_module;

  //cpu_3_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_3_jtag_debug_module_any_bursting_master_saved_grant = 0;

  //cpu_3_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_3_jtag_debug_module_arb_share_counter_next_value = cpu_3_jtag_debug_module_firsttransfer ? (cpu_3_jtag_debug_module_arb_share_set_values - 1) : |cpu_3_jtag_debug_module_arb_share_counter ? (cpu_3_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_3_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_3_jtag_debug_module_allgrants = (|cpu_3_jtag_debug_module_grant_vector) |
    (|cpu_3_jtag_debug_module_grant_vector) |
    (|cpu_3_jtag_debug_module_grant_vector) |
    (|cpu_3_jtag_debug_module_grant_vector);

  //cpu_3_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_3_jtag_debug_module_end_xfer = ~(cpu_3_jtag_debug_module_waits_for_read | cpu_3_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_3_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_3_jtag_debug_module = cpu_3_jtag_debug_module_end_xfer & (~cpu_3_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_3_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_3_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_3_jtag_debug_module & cpu_3_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_3_jtag_debug_module & ~cpu_3_jtag_debug_module_non_bursting_master_requests);

  //cpu_3_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_3_jtag_debug_module_arb_counter_enable)
          cpu_3_jtag_debug_module_arb_share_counter <= cpu_3_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_3_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_3_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_3_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_3_jtag_debug_module & ~cpu_3_jtag_debug_module_non_bursting_master_requests))
          cpu_3_jtag_debug_module_slavearbiterlockenable <= |cpu_3_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_3/data_master cpu_3/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = cpu_3_jtag_debug_module_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_3_jtag_debug_module_slavearbiterlockenable2 = |cpu_3_jtag_debug_module_arb_share_counter_next_value;

  //cpu_3/data_master cpu_3/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = cpu_3_jtag_debug_module_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/instruction_master cpu_3/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock = cpu_3_jtag_debug_module_slavearbiterlockenable & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master cpu_3/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock2 = cpu_3_jtag_debug_module_slavearbiterlockenable2 & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master granted cpu_3/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_instruction_master_granted_slave_cpu_3_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_3_instruction_master_granted_slave_cpu_3_jtag_debug_module <= cpu_3_instruction_master_saved_grant_cpu_3_jtag_debug_module ? 1 : (cpu_3_jtag_debug_module_arbitration_holdoff_internal | ~cpu_3_instruction_master_requests_cpu_3_jtag_debug_module) ? 0 : last_cycle_cpu_3_instruction_master_granted_slave_cpu_3_jtag_debug_module;
    end


  //cpu_3_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_3_instruction_master_continuerequest = last_cycle_cpu_3_instruction_master_granted_slave_cpu_3_jtag_debug_module & cpu_3_instruction_master_requests_cpu_3_jtag_debug_module;

  //cpu_3_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_3_jtag_debug_module_any_continuerequest = cpu_3_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest;

  assign cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module = cpu_3_data_master_requests_cpu_3_jtag_debug_module & ~((cpu_3_data_master_read & ((cpu_3_data_master_latency_counter != 0) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_3_instruction_master_arbiterlock);
  //local readdatavalid cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module, which is an e_mux
  assign cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module = cpu_3_data_master_granted_cpu_3_jtag_debug_module & cpu_3_data_master_read & ~cpu_3_jtag_debug_module_waits_for_read;

  //cpu_3_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_3_jtag_debug_module_writedata = cpu_3_data_master_writedata;

  assign cpu_3_instruction_master_requests_cpu_3_jtag_debug_module = (({cpu_3_instruction_master_address_to_slave[24 : 11] , 11'b0} == 25'h2000) & (cpu_3_instruction_master_read)) & cpu_3_instruction_master_read;
  //cpu_3/data_master granted cpu_3/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_cpu_3_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_cpu_3_jtag_debug_module <= cpu_3_data_master_saved_grant_cpu_3_jtag_debug_module ? 1 : (cpu_3_jtag_debug_module_arbitration_holdoff_internal | ~cpu_3_data_master_requests_cpu_3_jtag_debug_module) ? 0 : last_cycle_cpu_3_data_master_granted_slave_cpu_3_jtag_debug_module;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = last_cycle_cpu_3_data_master_granted_slave_cpu_3_jtag_debug_module & cpu_3_data_master_requests_cpu_3_jtag_debug_module;

  assign cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module = cpu_3_instruction_master_requests_cpu_3_jtag_debug_module & ~((cpu_3_instruction_master_read & ((cpu_3_instruction_master_latency_counter != 0) | (|cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module, which is an e_mux
  assign cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module = cpu_3_instruction_master_granted_cpu_3_jtag_debug_module & cpu_3_instruction_master_read & ~cpu_3_jtag_debug_module_waits_for_read;

  //allow new arb cycle for cpu_3/jtag_debug_module, which is an e_assign
  assign cpu_3_jtag_debug_module_allow_new_arb_cycle = ~cpu_3_data_master_arbiterlock & ~cpu_3_instruction_master_arbiterlock;

  //cpu_3/instruction_master assignment into master qualified-requests vector for cpu_3/jtag_debug_module, which is an e_assign
  assign cpu_3_jtag_debug_module_master_qreq_vector[0] = cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module;

  //cpu_3/instruction_master grant cpu_3/jtag_debug_module, which is an e_assign
  assign cpu_3_instruction_master_granted_cpu_3_jtag_debug_module = cpu_3_jtag_debug_module_grant_vector[0];

  //cpu_3/instruction_master saved-grant cpu_3/jtag_debug_module, which is an e_assign
  assign cpu_3_instruction_master_saved_grant_cpu_3_jtag_debug_module = cpu_3_jtag_debug_module_arb_winner[0] && cpu_3_instruction_master_requests_cpu_3_jtag_debug_module;

  //cpu_3/data_master assignment into master qualified-requests vector for cpu_3/jtag_debug_module, which is an e_assign
  assign cpu_3_jtag_debug_module_master_qreq_vector[1] = cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module;

  //cpu_3/data_master grant cpu_3/jtag_debug_module, which is an e_assign
  assign cpu_3_data_master_granted_cpu_3_jtag_debug_module = cpu_3_jtag_debug_module_grant_vector[1];

  //cpu_3/data_master saved-grant cpu_3/jtag_debug_module, which is an e_assign
  assign cpu_3_data_master_saved_grant_cpu_3_jtag_debug_module = cpu_3_jtag_debug_module_arb_winner[1] && cpu_3_data_master_requests_cpu_3_jtag_debug_module;

  //cpu_3/jtag_debug_module chosen-master double-vector, which is an e_assign
  assign cpu_3_jtag_debug_module_chosen_master_double_vector = {cpu_3_jtag_debug_module_master_qreq_vector, cpu_3_jtag_debug_module_master_qreq_vector} & ({~cpu_3_jtag_debug_module_master_qreq_vector, ~cpu_3_jtag_debug_module_master_qreq_vector} + cpu_3_jtag_debug_module_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_3_jtag_debug_module_arb_winner = (cpu_3_jtag_debug_module_allow_new_arb_cycle & | cpu_3_jtag_debug_module_grant_vector) ? cpu_3_jtag_debug_module_grant_vector : cpu_3_jtag_debug_module_saved_chosen_master_vector;

  //saved cpu_3_jtag_debug_module_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_jtag_debug_module_saved_chosen_master_vector <= 0;
      else if (cpu_3_jtag_debug_module_allow_new_arb_cycle)
          cpu_3_jtag_debug_module_saved_chosen_master_vector <= |cpu_3_jtag_debug_module_grant_vector ? cpu_3_jtag_debug_module_grant_vector : cpu_3_jtag_debug_module_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_3_jtag_debug_module_grant_vector = {(cpu_3_jtag_debug_module_chosen_master_double_vector[1] | cpu_3_jtag_debug_module_chosen_master_double_vector[3]),
    (cpu_3_jtag_debug_module_chosen_master_double_vector[0] | cpu_3_jtag_debug_module_chosen_master_double_vector[2])};

  //cpu_3/jtag_debug_module chosen master rotated left, which is an e_assign
  assign cpu_3_jtag_debug_module_chosen_master_rot_left = (cpu_3_jtag_debug_module_arb_winner << 1) ? (cpu_3_jtag_debug_module_arb_winner << 1) : 1;

  //cpu_3/jtag_debug_module's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_jtag_debug_module_arb_addend <= 1;
      else if (|cpu_3_jtag_debug_module_grant_vector)
          cpu_3_jtag_debug_module_arb_addend <= cpu_3_jtag_debug_module_end_xfer? cpu_3_jtag_debug_module_chosen_master_rot_left : cpu_3_jtag_debug_module_grant_vector;
    end


  assign cpu_3_jtag_debug_module_begintransfer = cpu_3_jtag_debug_module_begins_xfer;
  //assign cpu_3_jtag_debug_module_resetrequest_from_sa = cpu_3_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_3_jtag_debug_module_resetrequest_from_sa = cpu_3_jtag_debug_module_resetrequest;

  assign cpu_3_jtag_debug_module_chipselect = cpu_3_data_master_granted_cpu_3_jtag_debug_module | cpu_3_instruction_master_granted_cpu_3_jtag_debug_module;
  //cpu_3_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_3_jtag_debug_module_firsttransfer = cpu_3_jtag_debug_module_begins_xfer ? cpu_3_jtag_debug_module_unreg_firsttransfer : cpu_3_jtag_debug_module_reg_firsttransfer;

  //cpu_3_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_3_jtag_debug_module_unreg_firsttransfer = ~(cpu_3_jtag_debug_module_slavearbiterlockenable & cpu_3_jtag_debug_module_any_continuerequest);

  //cpu_3_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_3_jtag_debug_module_begins_xfer)
          cpu_3_jtag_debug_module_reg_firsttransfer <= cpu_3_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_3_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_3_jtag_debug_module_beginbursttransfer_internal = cpu_3_jtag_debug_module_begins_xfer;

  //cpu_3_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_3_jtag_debug_module_arbitration_holdoff_internal = cpu_3_jtag_debug_module_begins_xfer & cpu_3_jtag_debug_module_firsttransfer;

  //cpu_3_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_3_jtag_debug_module_write = cpu_3_data_master_granted_cpu_3_jtag_debug_module & cpu_3_data_master_write;

  assign shifted_address_to_cpu_3_jtag_debug_module_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  //cpu_3_jtag_debug_module_address mux, which is an e_mux
  assign cpu_3_jtag_debug_module_address = (cpu_3_data_master_granted_cpu_3_jtag_debug_module)? (shifted_address_to_cpu_3_jtag_debug_module_from_cpu_3_data_master >> 2) :
    (shifted_address_to_cpu_3_jtag_debug_module_from_cpu_3_instruction_master >> 2);

  assign shifted_address_to_cpu_3_jtag_debug_module_from_cpu_3_instruction_master = cpu_3_instruction_master_address_to_slave;
  //d1_cpu_3_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_3_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_3_jtag_debug_module_end_xfer <= cpu_3_jtag_debug_module_end_xfer;
    end


  //cpu_3_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_3_jtag_debug_module_waits_for_read = cpu_3_jtag_debug_module_in_a_read_cycle & cpu_3_jtag_debug_module_begins_xfer;

  //cpu_3_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_3_jtag_debug_module_in_a_read_cycle = (cpu_3_data_master_granted_cpu_3_jtag_debug_module & cpu_3_data_master_read) | (cpu_3_instruction_master_granted_cpu_3_jtag_debug_module & cpu_3_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_3_jtag_debug_module_in_a_read_cycle;

  //cpu_3_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_3_jtag_debug_module_waits_for_write = cpu_3_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_3_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_3_jtag_debug_module_in_a_write_cycle = cpu_3_data_master_granted_cpu_3_jtag_debug_module & cpu_3_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_3_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_3_jtag_debug_module_counter = 0;
  //cpu_3_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_3_jtag_debug_module_byteenable = (cpu_3_data_master_granted_cpu_3_jtag_debug_module)? cpu_3_data_master_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_3_jtag_debug_module_debugaccess = (cpu_3_data_master_granted_cpu_3_jtag_debug_module)? cpu_3_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_3/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_3_data_master_granted_cpu_3_jtag_debug_module + cpu_3_instruction_master_granted_cpu_3_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_3_data_master_saved_grant_cpu_3_jtag_debug_module + cpu_3_instruction_master_saved_grant_cpu_3_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_3_custom_instruction_master_arbitrator (
                                                    // inputs:
                                                     clk,
                                                     cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa,
                                                     cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa,
                                                     cpu_3_custom_instruction_master_multi_start,
                                                     reset_n,

                                                    // outputs:
                                                     cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select,
                                                     cpu_3_custom_instruction_master_multi_done,
                                                     cpu_3_custom_instruction_master_multi_result,
                                                     cpu_3_custom_instruction_master_reset_n,
                                                     cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1
                                                  )
;

  output           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select;
  output           cpu_3_custom_instruction_master_multi_done;
  output  [ 31: 0] cpu_3_custom_instruction_master_multi_result;
  output           cpu_3_custom_instruction_master_reset_n;
  output           cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1;
  input            clk;
  input            cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  input   [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  input            cpu_3_custom_instruction_master_multi_start;
  input            reset_n;

  wire             cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select;
  wire             cpu_3_custom_instruction_master_multi_done;
  wire    [ 31: 0] cpu_3_custom_instruction_master_multi_result;
  wire             cpu_3_custom_instruction_master_reset_n;
  wire             cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1;
  assign cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select = 1'b1;
  assign cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1 = cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select & cpu_3_custom_instruction_master_multi_start;
  //cpu_3_custom_instruction_master_multi_result mux, which is an e_mux
  assign cpu_3_custom_instruction_master_multi_result = {32 {cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select}} & cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;

  //multi_done mux, which is an e_mux
  assign cpu_3_custom_instruction_master_multi_done = {1 {cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select}} & cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;

  //cpu_3_custom_instruction_master_reset_n local reset_n, which is an e_assign
  assign cpu_3_custom_instruction_master_reset_n = reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_3_data_master_arbitrator (
                                      // inputs:
                                       clk,
                                       cpu_3_data_master_address,
                                       cpu_3_data_master_byteenable,
                                       cpu_3_data_master_byteenable_nios_system_clock_11_in,
                                       cpu_3_data_master_byteenable_nios_system_clock_7_in,
                                       cpu_3_data_master_byteenable_sram_0_avalon_sram_slave,
                                       cpu_3_data_master_granted_cpu_3_jtag_debug_module,
                                       cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave,
                                       cpu_3_data_master_granted_keys_s1,
                                       cpu_3_data_master_granted_mailbox_0_s1,
                                       cpu_3_data_master_granted_mailbox_1_s1,
                                       cpu_3_data_master_granted_mailbox_2_s1,
                                       cpu_3_data_master_granted_mailbox_3_s1,
                                       cpu_3_data_master_granted_nios_system_clock_11_in,
                                       cpu_3_data_master_granted_nios_system_clock_7_in,
                                       cpu_3_data_master_granted_onchip_memory2_0_s1,
                                       cpu_3_data_master_granted_onchip_memory2_1_s1,
                                       cpu_3_data_master_granted_onchip_memory2_2_s1,
                                       cpu_3_data_master_granted_onchip_memory2_3_s1,
                                       cpu_3_data_master_granted_performance_counter_0_control_slave,
                                       cpu_3_data_master_granted_sram_0_avalon_sram_slave,
                                       cpu_3_data_master_granted_sysid_control_slave,
                                       cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module,
                                       cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave,
                                       cpu_3_data_master_qualified_request_keys_s1,
                                       cpu_3_data_master_qualified_request_mailbox_0_s1,
                                       cpu_3_data_master_qualified_request_mailbox_1_s1,
                                       cpu_3_data_master_qualified_request_mailbox_2_s1,
                                       cpu_3_data_master_qualified_request_mailbox_3_s1,
                                       cpu_3_data_master_qualified_request_nios_system_clock_11_in,
                                       cpu_3_data_master_qualified_request_nios_system_clock_7_in,
                                       cpu_3_data_master_qualified_request_onchip_memory2_0_s1,
                                       cpu_3_data_master_qualified_request_onchip_memory2_1_s1,
                                       cpu_3_data_master_qualified_request_onchip_memory2_2_s1,
                                       cpu_3_data_master_qualified_request_onchip_memory2_3_s1,
                                       cpu_3_data_master_qualified_request_performance_counter_0_control_slave,
                                       cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave,
                                       cpu_3_data_master_qualified_request_sysid_control_slave,
                                       cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_3_data_master_read,
                                       cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module,
                                       cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave,
                                       cpu_3_data_master_read_data_valid_keys_s1,
                                       cpu_3_data_master_read_data_valid_mailbox_0_s1,
                                       cpu_3_data_master_read_data_valid_mailbox_1_s1,
                                       cpu_3_data_master_read_data_valid_mailbox_2_s1,
                                       cpu_3_data_master_read_data_valid_mailbox_3_s1,
                                       cpu_3_data_master_read_data_valid_nios_system_clock_11_in,
                                       cpu_3_data_master_read_data_valid_nios_system_clock_7_in,
                                       cpu_3_data_master_read_data_valid_onchip_memory2_0_s1,
                                       cpu_3_data_master_read_data_valid_onchip_memory2_1_s1,
                                       cpu_3_data_master_read_data_valid_onchip_memory2_2_s1,
                                       cpu_3_data_master_read_data_valid_onchip_memory2_3_s1,
                                       cpu_3_data_master_read_data_valid_performance_counter_0_control_slave,
                                       cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave,
                                       cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                       cpu_3_data_master_read_data_valid_sysid_control_slave,
                                       cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_3_data_master_requests_cpu_3_jtag_debug_module,
                                       cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave,
                                       cpu_3_data_master_requests_keys_s1,
                                       cpu_3_data_master_requests_mailbox_0_s1,
                                       cpu_3_data_master_requests_mailbox_1_s1,
                                       cpu_3_data_master_requests_mailbox_2_s1,
                                       cpu_3_data_master_requests_mailbox_3_s1,
                                       cpu_3_data_master_requests_nios_system_clock_11_in,
                                       cpu_3_data_master_requests_nios_system_clock_7_in,
                                       cpu_3_data_master_requests_onchip_memory2_0_s1,
                                       cpu_3_data_master_requests_onchip_memory2_1_s1,
                                       cpu_3_data_master_requests_onchip_memory2_2_s1,
                                       cpu_3_data_master_requests_onchip_memory2_3_s1,
                                       cpu_3_data_master_requests_performance_counter_0_control_slave,
                                       cpu_3_data_master_requests_sram_0_avalon_sram_slave,
                                       cpu_3_data_master_requests_sysid_control_slave,
                                       cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave,
                                       cpu_3_data_master_write,
                                       cpu_3_data_master_writedata,
                                       cpu_3_jtag_debug_module_readdata_from_sa,
                                       d1_cpu_3_jtag_debug_module_end_xfer,
                                       d1_jtag_uart_3_avalon_jtag_slave_end_xfer,
                                       d1_keys_s1_end_xfer,
                                       d1_mailbox_0_s1_end_xfer,
                                       d1_mailbox_1_s1_end_xfer,
                                       d1_mailbox_2_s1_end_xfer,
                                       d1_mailbox_3_s1_end_xfer,
                                       d1_nios_system_clock_11_in_end_xfer,
                                       d1_nios_system_clock_7_in_end_xfer,
                                       d1_onchip_memory2_0_s1_end_xfer,
                                       d1_onchip_memory2_1_s1_end_xfer,
                                       d1_onchip_memory2_2_s1_end_xfer,
                                       d1_onchip_memory2_3_s1_end_xfer,
                                       d1_performance_counter_0_control_slave_end_xfer,
                                       d1_sram_0_avalon_sram_slave_end_xfer,
                                       d1_sysid_control_slave_end_xfer,
                                       d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer,
                                       jtag_uart_3_avalon_jtag_slave_irq_from_sa,
                                       jtag_uart_3_avalon_jtag_slave_readdata_from_sa,
                                       jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa,
                                       keys_s1_readdata_from_sa,
                                       mailbox_0_s1_readdata_from_sa,
                                       mailbox_1_s1_readdata_from_sa,
                                       mailbox_2_s1_readdata_from_sa,
                                       mailbox_3_s1_readdata_from_sa,
                                       nios_system_clock_11_in_readdata_from_sa,
                                       nios_system_clock_11_in_waitrequest_from_sa,
                                       nios_system_clock_7_in_readdata_from_sa,
                                       nios_system_clock_7_in_waitrequest_from_sa,
                                       onchip_memory2_0_s1_readdata_from_sa,
                                       onchip_memory2_1_s1_readdata_from_sa,
                                       onchip_memory2_2_s1_readdata_from_sa,
                                       onchip_memory2_3_s1_readdata_from_sa,
                                       performance_counter_0_control_slave_readdata_from_sa,
                                       reset_n,
                                       sram_0_avalon_sram_slave_readdata_from_sa,
                                       sysid_control_slave_readdata_from_sa,
                                       video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa,

                                      // outputs:
                                       cpu_3_data_master_address_to_slave,
                                       cpu_3_data_master_dbs_address,
                                       cpu_3_data_master_dbs_write_16,
                                       cpu_3_data_master_dbs_write_8,
                                       cpu_3_data_master_irq,
                                       cpu_3_data_master_latency_counter,
                                       cpu_3_data_master_readdata,
                                       cpu_3_data_master_readdatavalid,
                                       cpu_3_data_master_waitrequest
                                    )
;

  output  [ 24: 0] cpu_3_data_master_address_to_slave;
  output  [  1: 0] cpu_3_data_master_dbs_address;
  output  [ 15: 0] cpu_3_data_master_dbs_write_16;
  output  [  7: 0] cpu_3_data_master_dbs_write_8;
  output  [ 31: 0] cpu_3_data_master_irq;
  output           cpu_3_data_master_latency_counter;
  output  [ 31: 0] cpu_3_data_master_readdata;
  output           cpu_3_data_master_readdatavalid;
  output           cpu_3_data_master_waitrequest;
  input            clk;
  input   [ 24: 0] cpu_3_data_master_address;
  input   [  3: 0] cpu_3_data_master_byteenable;
  input            cpu_3_data_master_byteenable_nios_system_clock_11_in;
  input   [  1: 0] cpu_3_data_master_byteenable_nios_system_clock_7_in;
  input   [  1: 0] cpu_3_data_master_byteenable_sram_0_avalon_sram_slave;
  input            cpu_3_data_master_granted_cpu_3_jtag_debug_module;
  input            cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave;
  input            cpu_3_data_master_granted_keys_s1;
  input            cpu_3_data_master_granted_mailbox_0_s1;
  input            cpu_3_data_master_granted_mailbox_1_s1;
  input            cpu_3_data_master_granted_mailbox_2_s1;
  input            cpu_3_data_master_granted_mailbox_3_s1;
  input            cpu_3_data_master_granted_nios_system_clock_11_in;
  input            cpu_3_data_master_granted_nios_system_clock_7_in;
  input            cpu_3_data_master_granted_onchip_memory2_0_s1;
  input            cpu_3_data_master_granted_onchip_memory2_1_s1;
  input            cpu_3_data_master_granted_onchip_memory2_2_s1;
  input            cpu_3_data_master_granted_onchip_memory2_3_s1;
  input            cpu_3_data_master_granted_performance_counter_0_control_slave;
  input            cpu_3_data_master_granted_sram_0_avalon_sram_slave;
  input            cpu_3_data_master_granted_sysid_control_slave;
  input            cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module;
  input            cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave;
  input            cpu_3_data_master_qualified_request_keys_s1;
  input            cpu_3_data_master_qualified_request_mailbox_0_s1;
  input            cpu_3_data_master_qualified_request_mailbox_1_s1;
  input            cpu_3_data_master_qualified_request_mailbox_2_s1;
  input            cpu_3_data_master_qualified_request_mailbox_3_s1;
  input            cpu_3_data_master_qualified_request_nios_system_clock_11_in;
  input            cpu_3_data_master_qualified_request_nios_system_clock_7_in;
  input            cpu_3_data_master_qualified_request_onchip_memory2_0_s1;
  input            cpu_3_data_master_qualified_request_onchip_memory2_1_s1;
  input            cpu_3_data_master_qualified_request_onchip_memory2_2_s1;
  input            cpu_3_data_master_qualified_request_onchip_memory2_3_s1;
  input            cpu_3_data_master_qualified_request_performance_counter_0_control_slave;
  input            cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave;
  input            cpu_3_data_master_qualified_request_sysid_control_slave;
  input            cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module;
  input            cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave;
  input            cpu_3_data_master_read_data_valid_keys_s1;
  input            cpu_3_data_master_read_data_valid_mailbox_0_s1;
  input            cpu_3_data_master_read_data_valid_mailbox_1_s1;
  input            cpu_3_data_master_read_data_valid_mailbox_2_s1;
  input            cpu_3_data_master_read_data_valid_mailbox_3_s1;
  input            cpu_3_data_master_read_data_valid_nios_system_clock_11_in;
  input            cpu_3_data_master_read_data_valid_nios_system_clock_7_in;
  input            cpu_3_data_master_read_data_valid_onchip_memory2_0_s1;
  input            cpu_3_data_master_read_data_valid_onchip_memory2_1_s1;
  input            cpu_3_data_master_read_data_valid_onchip_memory2_2_s1;
  input            cpu_3_data_master_read_data_valid_onchip_memory2_3_s1;
  input            cpu_3_data_master_read_data_valid_performance_counter_0_control_slave;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_read_data_valid_sysid_control_slave;
  input            cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_3_data_master_requests_cpu_3_jtag_debug_module;
  input            cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave;
  input            cpu_3_data_master_requests_keys_s1;
  input            cpu_3_data_master_requests_mailbox_0_s1;
  input            cpu_3_data_master_requests_mailbox_1_s1;
  input            cpu_3_data_master_requests_mailbox_2_s1;
  input            cpu_3_data_master_requests_mailbox_3_s1;
  input            cpu_3_data_master_requests_nios_system_clock_11_in;
  input            cpu_3_data_master_requests_nios_system_clock_7_in;
  input            cpu_3_data_master_requests_onchip_memory2_0_s1;
  input            cpu_3_data_master_requests_onchip_memory2_1_s1;
  input            cpu_3_data_master_requests_onchip_memory2_2_s1;
  input            cpu_3_data_master_requests_onchip_memory2_3_s1;
  input            cpu_3_data_master_requests_performance_counter_0_control_slave;
  input            cpu_3_data_master_requests_sram_0_avalon_sram_slave;
  input            cpu_3_data_master_requests_sysid_control_slave;
  input            cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 31: 0] cpu_3_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_3_jtag_debug_module_end_xfer;
  input            d1_jtag_uart_3_avalon_jtag_slave_end_xfer;
  input            d1_keys_s1_end_xfer;
  input            d1_mailbox_0_s1_end_xfer;
  input            d1_mailbox_1_s1_end_xfer;
  input            d1_mailbox_2_s1_end_xfer;
  input            d1_mailbox_3_s1_end_xfer;
  input            d1_nios_system_clock_11_in_end_xfer;
  input            d1_nios_system_clock_7_in_end_xfer;
  input            d1_onchip_memory2_0_s1_end_xfer;
  input            d1_onchip_memory2_1_s1_end_xfer;
  input            d1_onchip_memory2_2_s1_end_xfer;
  input            d1_onchip_memory2_3_s1_end_xfer;
  input            d1_performance_counter_0_control_slave_end_xfer;
  input            d1_sram_0_avalon_sram_slave_end_xfer;
  input            d1_sysid_control_slave_end_xfer;
  input            d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer;
  input            jtag_uart_3_avalon_jtag_slave_irq_from_sa;
  input   [ 31: 0] jtag_uart_3_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa;
  input   [ 31: 0] keys_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_0_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_1_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_2_s1_readdata_from_sa;
  input   [ 31: 0] mailbox_3_s1_readdata_from_sa;
  input   [  7: 0] nios_system_clock_11_in_readdata_from_sa;
  input            nios_system_clock_11_in_waitrequest_from_sa;
  input   [ 15: 0] nios_system_clock_7_in_readdata_from_sa;
  input            nios_system_clock_7_in_waitrequest_from_sa;
  input   [ 31: 0] onchip_memory2_0_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_1_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_2_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_3_s1_readdata_from_sa;
  input   [ 31: 0] performance_counter_0_control_slave_readdata_from_sa;
  input            reset_n;
  input   [ 15: 0] sram_0_avalon_sram_slave_readdata_from_sa;
  input   [ 31: 0] sysid_control_slave_readdata_from_sa;
  input   [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] cpu_3_data_master_address_last_time;
  wire    [ 24: 0] cpu_3_data_master_address_to_slave;
  reg     [  3: 0] cpu_3_data_master_byteenable_last_time;
  reg     [  1: 0] cpu_3_data_master_dbs_address;
  wire    [  1: 0] cpu_3_data_master_dbs_increment;
  reg     [  1: 0] cpu_3_data_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_3_data_master_dbs_rdv_counter_inc;
  wire    [ 15: 0] cpu_3_data_master_dbs_write_16;
  wire    [  7: 0] cpu_3_data_master_dbs_write_8;
  wire    [ 31: 0] cpu_3_data_master_irq;
  wire             cpu_3_data_master_is_granted_some_slave;
  reg              cpu_3_data_master_latency_counter;
  wire    [  1: 0] cpu_3_data_master_next_dbs_rdv_counter;
  reg              cpu_3_data_master_read_but_no_slave_selected;
  reg              cpu_3_data_master_read_last_time;
  wire    [ 31: 0] cpu_3_data_master_readdata;
  wire             cpu_3_data_master_readdatavalid;
  wire             cpu_3_data_master_run;
  wire             cpu_3_data_master_waitrequest;
  reg              cpu_3_data_master_write_last_time;
  reg     [ 31: 0] cpu_3_data_master_writedata_last_time;
  reg     [ 15: 0] dbs_16_reg_segment_0;
  reg     [  7: 0] dbs_8_reg_segment_0;
  reg     [  7: 0] dbs_8_reg_segment_1;
  reg     [  7: 0] dbs_8_reg_segment_2;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire             p1_cpu_3_data_master_latency_counter;
  wire    [ 15: 0] p1_dbs_16_reg_segment_0;
  wire    [  7: 0] p1_dbs_8_reg_segment_0;
  wire    [  7: 0] p1_dbs_8_reg_segment_1;
  wire    [  7: 0] p1_dbs_8_reg_segment_2;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_3_data_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  wire             r_3;
  wire             r_4;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module | ~cpu_3_data_master_requests_cpu_3_jtag_debug_module) & (cpu_3_data_master_granted_cpu_3_jtag_debug_module | ~cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module) & ((~cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module | ~cpu_3_data_master_read | (1 & ~d1_cpu_3_jtag_debug_module_end_xfer & cpu_3_data_master_read))) & ((~cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module | ~cpu_3_data_master_write | (1 & cpu_3_data_master_write))) & 1 & (cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave | ~cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave) & ((~cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & ~jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa & (cpu_3_data_master_read | cpu_3_data_master_write)))) & ((~cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & ~jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa & (cpu_3_data_master_read | cpu_3_data_master_write)))) & 1 & (cpu_3_data_master_qualified_request_keys_s1 | ~cpu_3_data_master_requests_keys_s1) & (cpu_3_data_master_granted_keys_s1 | ~cpu_3_data_master_qualified_request_keys_s1) & ((~cpu_3_data_master_qualified_request_keys_s1 | ~cpu_3_data_master_read | (1 & ~d1_keys_s1_end_xfer & cpu_3_data_master_read))) & ((~cpu_3_data_master_qualified_request_keys_s1 | ~cpu_3_data_master_write | (1 & cpu_3_data_master_write))) & 1 & (cpu_3_data_master_qualified_request_mailbox_0_s1 | ~cpu_3_data_master_requests_mailbox_0_s1) & (cpu_3_data_master_granted_mailbox_0_s1 | ~cpu_3_data_master_qualified_request_mailbox_0_s1) & ((~cpu_3_data_master_qualified_request_mailbox_0_s1 | ~cpu_3_data_master_read | (1 & ~d1_mailbox_0_s1_end_xfer & cpu_3_data_master_read))) & ((~cpu_3_data_master_qualified_request_mailbox_0_s1 | ~cpu_3_data_master_write | (1 & cpu_3_data_master_write)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_3_data_master_run = r_0 & r_1 & r_2 & r_3 & r_4;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_3_data_master_qualified_request_mailbox_1_s1 | ~cpu_3_data_master_requests_mailbox_1_s1) & (cpu_3_data_master_granted_mailbox_1_s1 | ~cpu_3_data_master_qualified_request_mailbox_1_s1) & ((~cpu_3_data_master_qualified_request_mailbox_1_s1 | ~cpu_3_data_master_read | (1 & ~d1_mailbox_1_s1_end_xfer & cpu_3_data_master_read))) & ((~cpu_3_data_master_qualified_request_mailbox_1_s1 | ~cpu_3_data_master_write | (1 & cpu_3_data_master_write))) & 1 & (cpu_3_data_master_qualified_request_mailbox_2_s1 | ~cpu_3_data_master_requests_mailbox_2_s1) & (cpu_3_data_master_granted_mailbox_2_s1 | ~cpu_3_data_master_qualified_request_mailbox_2_s1) & ((~cpu_3_data_master_qualified_request_mailbox_2_s1 | ~cpu_3_data_master_read | (1 & ~d1_mailbox_2_s1_end_xfer & cpu_3_data_master_read))) & ((~cpu_3_data_master_qualified_request_mailbox_2_s1 | ~cpu_3_data_master_write | (1 & cpu_3_data_master_write))) & 1 & (cpu_3_data_master_qualified_request_mailbox_3_s1 | ~cpu_3_data_master_requests_mailbox_3_s1) & (cpu_3_data_master_granted_mailbox_3_s1 | ~cpu_3_data_master_qualified_request_mailbox_3_s1) & ((~cpu_3_data_master_qualified_request_mailbox_3_s1 | ~cpu_3_data_master_read | (1 & ~d1_mailbox_3_s1_end_xfer & cpu_3_data_master_read))) & ((~cpu_3_data_master_qualified_request_mailbox_3_s1 | ~cpu_3_data_master_write | (1 & cpu_3_data_master_write))) & 1 & ((cpu_3_data_master_qualified_request_nios_system_clock_11_in | ((cpu_3_data_master_write & !cpu_3_data_master_byteenable_nios_system_clock_11_in & cpu_3_data_master_dbs_address[1] & cpu_3_data_master_dbs_address[0])) | ~cpu_3_data_master_requests_nios_system_clock_11_in)) & ((~cpu_3_data_master_qualified_request_nios_system_clock_11_in | ~cpu_3_data_master_read | (1 & ~nios_system_clock_11_in_waitrequest_from_sa & (cpu_3_data_master_dbs_address[1] & cpu_3_data_master_dbs_address[0]) & cpu_3_data_master_read))) & ((~cpu_3_data_master_qualified_request_nios_system_clock_11_in | ~cpu_3_data_master_write | (1 & ~nios_system_clock_11_in_waitrequest_from_sa & (cpu_3_data_master_dbs_address[1] & cpu_3_data_master_dbs_address[0]) & cpu_3_data_master_write)));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_3_data_master_qualified_request_nios_system_clock_7_in | (cpu_3_data_master_write & !cpu_3_data_master_byteenable_nios_system_clock_7_in & cpu_3_data_master_dbs_address[1]) | ~cpu_3_data_master_requests_nios_system_clock_7_in) & ((~cpu_3_data_master_qualified_request_nios_system_clock_7_in | ~cpu_3_data_master_read | (1 & ~nios_system_clock_7_in_waitrequest_from_sa & (cpu_3_data_master_dbs_address[1]) & cpu_3_data_master_read))) & ((~cpu_3_data_master_qualified_request_nios_system_clock_7_in | ~cpu_3_data_master_write | (1 & ~nios_system_clock_7_in_waitrequest_from_sa & (cpu_3_data_master_dbs_address[1]) & cpu_3_data_master_write))) & 1 & (cpu_3_data_master_qualified_request_onchip_memory2_0_s1 | ~cpu_3_data_master_requests_onchip_memory2_0_s1) & (cpu_3_data_master_granted_onchip_memory2_0_s1 | ~cpu_3_data_master_qualified_request_onchip_memory2_0_s1) & ((~cpu_3_data_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write)))) & ((~cpu_3_data_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write)))) & 1 & (cpu_3_data_master_qualified_request_onchip_memory2_1_s1 | ~cpu_3_data_master_requests_onchip_memory2_1_s1) & (cpu_3_data_master_granted_onchip_memory2_1_s1 | ~cpu_3_data_master_qualified_request_onchip_memory2_1_s1) & ((~cpu_3_data_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write)))) & ((~cpu_3_data_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write)))) & 1 & (cpu_3_data_master_qualified_request_onchip_memory2_2_s1 | ~cpu_3_data_master_requests_onchip_memory2_2_s1) & (cpu_3_data_master_granted_onchip_memory2_2_s1 | ~cpu_3_data_master_qualified_request_onchip_memory2_2_s1) & ((~cpu_3_data_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write)))) & ((~cpu_3_data_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write))));

  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (cpu_3_data_master_qualified_request_onchip_memory2_3_s1 | ~cpu_3_data_master_requests_onchip_memory2_3_s1) & (cpu_3_data_master_granted_onchip_memory2_3_s1 | ~cpu_3_data_master_qualified_request_onchip_memory2_3_s1) & ((~cpu_3_data_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write)))) & ((~cpu_3_data_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write)))) & 1 & (cpu_3_data_master_qualified_request_performance_counter_0_control_slave | ~cpu_3_data_master_requests_performance_counter_0_control_slave) & (cpu_3_data_master_granted_performance_counter_0_control_slave | ~cpu_3_data_master_qualified_request_performance_counter_0_control_slave) & ((~cpu_3_data_master_qualified_request_performance_counter_0_control_slave | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write)))) & ((~cpu_3_data_master_qualified_request_performance_counter_0_control_slave | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write)))) & 1 & (cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave | (cpu_3_data_master_write & !cpu_3_data_master_byteenable_sram_0_avalon_sram_slave & cpu_3_data_master_dbs_address[1]) | ~cpu_3_data_master_requests_sram_0_avalon_sram_slave) & (cpu_3_data_master_granted_sram_0_avalon_sram_slave | ~cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave) & ((~cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_3_data_master_read | (1 & (cpu_3_data_master_dbs_address[1]) & cpu_3_data_master_read))) & ((~cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_3_data_master_write | (1 & (cpu_3_data_master_dbs_address[1]) & cpu_3_data_master_write))) & 1 & (cpu_3_data_master_qualified_request_sysid_control_slave | ~cpu_3_data_master_requests_sysid_control_slave) & (cpu_3_data_master_granted_sysid_control_slave | ~cpu_3_data_master_qualified_request_sysid_control_slave) & ((~cpu_3_data_master_qualified_request_sysid_control_slave | ~cpu_3_data_master_read | (1 & ~d1_sysid_control_slave_end_xfer & cpu_3_data_master_read)));

  //r_4 master_run cascaded wait assignment, which is an e_assign
  assign r_4 = ((~cpu_3_data_master_qualified_request_sysid_control_slave | ~cpu_3_data_master_write | (1 & cpu_3_data_master_write))) & 1 & (cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) & (cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave | ~cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave) & ((~cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write)))) & ((~cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | ~(cpu_3_data_master_read | cpu_3_data_master_write) | (1 & (cpu_3_data_master_read | cpu_3_data_master_write))));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_3_data_master_address_to_slave = cpu_3_data_master_address[24 : 0];

  //cpu_3_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_read_but_no_slave_selected <= 0;
      else 
        cpu_3_data_master_read_but_no_slave_selected <= cpu_3_data_master_read & cpu_3_data_master_run & ~cpu_3_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_3_data_master_is_granted_some_slave = cpu_3_data_master_granted_cpu_3_jtag_debug_module |
    cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave |
    cpu_3_data_master_granted_keys_s1 |
    cpu_3_data_master_granted_mailbox_0_s1 |
    cpu_3_data_master_granted_mailbox_1_s1 |
    cpu_3_data_master_granted_mailbox_2_s1 |
    cpu_3_data_master_granted_mailbox_3_s1 |
    cpu_3_data_master_granted_nios_system_clock_11_in |
    cpu_3_data_master_granted_nios_system_clock_7_in |
    cpu_3_data_master_granted_onchip_memory2_0_s1 |
    cpu_3_data_master_granted_onchip_memory2_1_s1 |
    cpu_3_data_master_granted_onchip_memory2_2_s1 |
    cpu_3_data_master_granted_onchip_memory2_3_s1 |
    cpu_3_data_master_granted_performance_counter_0_control_slave |
    cpu_3_data_master_granted_sram_0_avalon_sram_slave |
    cpu_3_data_master_granted_sysid_control_slave |
    cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_3_data_master_readdatavalid = cpu_3_data_master_read_data_valid_onchip_memory2_0_s1 |
    cpu_3_data_master_read_data_valid_onchip_memory2_1_s1 |
    cpu_3_data_master_read_data_valid_onchip_memory2_2_s1 |
    cpu_3_data_master_read_data_valid_onchip_memory2_3_s1 |
    cpu_3_data_master_read_data_valid_performance_counter_0_control_slave |
    (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave & dbs_rdv_counter_overflow) |
    cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_3_data_master_readdatavalid = cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_data_valid_keys_s1 |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_data_valid_mailbox_0_s1 |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_data_valid_mailbox_1_s1 |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_data_valid_mailbox_2_s1 |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_data_valid_mailbox_3_s1 |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    (cpu_3_data_master_read_data_valid_nios_system_clock_11_in & dbs_counter_overflow) |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    (cpu_3_data_master_read_data_valid_nios_system_clock_7_in & dbs_counter_overflow) |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid |
    cpu_3_data_master_read_data_valid_sysid_control_slave |
    cpu_3_data_master_read_but_no_slave_selected |
    pre_flush_cpu_3_data_master_readdatavalid;

  //cpu_3/data_master readdata mux, which is an e_mux
  assign cpu_3_data_master_readdata = ({32 {~(cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module & cpu_3_data_master_read)}} | cpu_3_jtag_debug_module_readdata_from_sa) &
    ({32 {~(cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave & cpu_3_data_master_read)}} | jtag_uart_3_avalon_jtag_slave_readdata_from_sa) &
    ({32 {~(cpu_3_data_master_qualified_request_keys_s1 & cpu_3_data_master_read)}} | keys_s1_readdata_from_sa) &
    ({32 {~(cpu_3_data_master_qualified_request_mailbox_0_s1 & cpu_3_data_master_read)}} | mailbox_0_s1_readdata_from_sa) &
    ({32 {~(cpu_3_data_master_qualified_request_mailbox_1_s1 & cpu_3_data_master_read)}} | mailbox_1_s1_readdata_from_sa) &
    ({32 {~(cpu_3_data_master_qualified_request_mailbox_2_s1 & cpu_3_data_master_read)}} | mailbox_2_s1_readdata_from_sa) &
    ({32 {~(cpu_3_data_master_qualified_request_mailbox_3_s1 & cpu_3_data_master_read)}} | mailbox_3_s1_readdata_from_sa) &
    ({32 {~(cpu_3_data_master_qualified_request_nios_system_clock_11_in & cpu_3_data_master_read)}} | {nios_system_clock_11_in_readdata_from_sa[7 : 0],
    dbs_8_reg_segment_2,
    dbs_8_reg_segment_1,
    dbs_8_reg_segment_0}) &
    ({32 {~(cpu_3_data_master_qualified_request_nios_system_clock_7_in & cpu_3_data_master_read)}} | {nios_system_clock_7_in_readdata_from_sa[15 : 0],
    dbs_16_reg_segment_0}) &
    ({32 {~cpu_3_data_master_read_data_valid_onchip_memory2_0_s1}} | onchip_memory2_0_s1_readdata_from_sa) &
    ({32 {~cpu_3_data_master_read_data_valid_onchip_memory2_1_s1}} | onchip_memory2_1_s1_readdata_from_sa) &
    ({32 {~cpu_3_data_master_read_data_valid_onchip_memory2_2_s1}} | onchip_memory2_2_s1_readdata_from_sa) &
    ({32 {~cpu_3_data_master_read_data_valid_onchip_memory2_3_s1}} | onchip_memory2_3_s1_readdata_from_sa) &
    ({32 {~cpu_3_data_master_read_data_valid_performance_counter_0_control_slave}} | performance_counter_0_control_slave_readdata_from_sa) &
    ({32 {~cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave}} | {sram_0_avalon_sram_slave_readdata_from_sa[15 : 0],
    dbs_latent_16_reg_segment_0}) &
    ({32 {~(cpu_3_data_master_qualified_request_sysid_control_slave & cpu_3_data_master_read)}} | sysid_control_slave_readdata_from_sa) &
    ({32 {~cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave}} | video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_3_data_master_waitrequest = ~cpu_3_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_latency_counter <= 0;
      else 
        cpu_3_data_master_latency_counter <= p1_cpu_3_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_3_data_master_latency_counter = ((cpu_3_data_master_run & cpu_3_data_master_read))? latency_load_value :
    (cpu_3_data_master_latency_counter)? cpu_3_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({1 {cpu_3_data_master_requests_onchip_memory2_0_s1}} & 1) |
    ({1 {cpu_3_data_master_requests_onchip_memory2_1_s1}} & 1) |
    ({1 {cpu_3_data_master_requests_onchip_memory2_2_s1}} & 1) |
    ({1 {cpu_3_data_master_requests_onchip_memory2_3_s1}} & 1) |
    ({1 {cpu_3_data_master_requests_performance_counter_0_control_slave}} & 1) |
    ({1 {cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave}} & 1);

  //irq assign, which is an e_assign
  assign cpu_3_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    jtag_uart_3_avalon_jtag_slave_irq_from_sa,
    1'b0};

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (((~0) & cpu_3_data_master_requests_nios_system_clock_11_in & cpu_3_data_master_write & !cpu_3_data_master_byteenable_nios_system_clock_11_in)) |
    (cpu_3_data_master_granted_nios_system_clock_11_in & cpu_3_data_master_read & 1 & 1 & ~nios_system_clock_11_in_waitrequest_from_sa) |
    (cpu_3_data_master_granted_nios_system_clock_11_in & cpu_3_data_master_write & 1 & 1 & ~nios_system_clock_11_in_waitrequest_from_sa) |
    (((~0) & cpu_3_data_master_requests_nios_system_clock_7_in & cpu_3_data_master_write & !cpu_3_data_master_byteenable_nios_system_clock_7_in)) |
    (cpu_3_data_master_granted_nios_system_clock_7_in & cpu_3_data_master_read & 1 & 1 & ~nios_system_clock_7_in_waitrequest_from_sa) |
    (cpu_3_data_master_granted_nios_system_clock_7_in & cpu_3_data_master_write & 1 & 1 & ~nios_system_clock_7_in_waitrequest_from_sa) |
    (((~0) & cpu_3_data_master_requests_sram_0_avalon_sram_slave & cpu_3_data_master_write & !cpu_3_data_master_byteenable_sram_0_avalon_sram_slave)) |
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave & cpu_3_data_master_read & 1 & 1) |
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave & cpu_3_data_master_write & 1 & 1);

  //input to dbs-8 stored 0, which is an e_mux
  assign p1_dbs_8_reg_segment_0 = nios_system_clock_11_in_readdata_from_sa;

  //dbs register for dbs-8 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_3_data_master_dbs_address[1 : 0]) == 0))
          dbs_8_reg_segment_0 <= p1_dbs_8_reg_segment_0;
    end


  //input to dbs-8 stored 1, which is an e_mux
  assign p1_dbs_8_reg_segment_1 = nios_system_clock_11_in_readdata_from_sa;

  //dbs register for dbs-8 segment 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_1 <= 0;
      else if (dbs_count_enable & ((cpu_3_data_master_dbs_address[1 : 0]) == 1))
          dbs_8_reg_segment_1 <= p1_dbs_8_reg_segment_1;
    end


  //input to dbs-8 stored 2, which is an e_mux
  assign p1_dbs_8_reg_segment_2 = nios_system_clock_11_in_readdata_from_sa;

  //dbs register for dbs-8 segment 2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_8_reg_segment_2 <= 0;
      else if (dbs_count_enable & ((cpu_3_data_master_dbs_address[1 : 0]) == 2))
          dbs_8_reg_segment_2 <= p1_dbs_8_reg_segment_2;
    end


  //mux write dbs 2, which is an e_mux
  assign cpu_3_data_master_dbs_write_8 = ((cpu_3_data_master_dbs_address[1 : 0] == 0))? cpu_3_data_master_writedata[7 : 0] :
    ((cpu_3_data_master_dbs_address[1 : 0] == 1))? cpu_3_data_master_writedata[15 : 8] :
    ((cpu_3_data_master_dbs_address[1 : 0] == 2))? cpu_3_data_master_writedata[23 : 16] :
    cpu_3_data_master_writedata[31 : 24];

  //dbs count increment, which is an e_mux
  assign cpu_3_data_master_dbs_increment = (cpu_3_data_master_requests_nios_system_clock_11_in)? 1 :
    (cpu_3_data_master_requests_nios_system_clock_7_in)? 2 :
    (cpu_3_data_master_requests_sram_0_avalon_sram_slave)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_3_data_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_3_data_master_dbs_address + cpu_3_data_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_3_data_master_dbs_address <= next_dbs_address;
    end


  //input to dbs-16 stored 0, which is an e_mux
  assign p1_dbs_16_reg_segment_0 = nios_system_clock_7_in_readdata_from_sa;

  //dbs register for dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_16_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_3_data_master_dbs_address[1]) == 0))
          dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
    end


  //mux write dbs 1, which is an e_mux
  assign cpu_3_data_master_dbs_write_16 = (cpu_3_data_master_dbs_address[1])? cpu_3_data_master_writedata[31 : 16] :
    (~(cpu_3_data_master_dbs_address[1]))? cpu_3_data_master_writedata[15 : 0] :
    (cpu_3_data_master_dbs_address[1])? cpu_3_data_master_writedata[31 : 16] :
    cpu_3_data_master_writedata[15 : 0];

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = sram_0_avalon_sram_slave_readdata_from_sa;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_3_data_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_3_data_master_next_dbs_rdv_counter = cpu_3_data_master_dbs_rdv_counter + cpu_3_data_master_dbs_rdv_counter_inc;

  //cpu_3_data_master_rdv_inc_mux, which is an e_mux
  assign cpu_3_data_master_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_3_data_master_dbs_rdv_counter <= cpu_3_data_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_3_data_master_dbs_rdv_counter[1] & ~cpu_3_data_master_next_dbs_rdv_counter[1];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_3_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_address_last_time <= 0;
      else 
        cpu_3_data_master_address_last_time <= cpu_3_data_master_address;
    end


  //cpu_3/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_3_data_master_waitrequest & (cpu_3_data_master_read | cpu_3_data_master_write);
    end


  //cpu_3_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_3_data_master_address != cpu_3_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_3_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_3_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_byteenable_last_time <= 0;
      else 
        cpu_3_data_master_byteenable_last_time <= cpu_3_data_master_byteenable;
    end


  //cpu_3_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_3_data_master_byteenable != cpu_3_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_3_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_3_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_read_last_time <= 0;
      else 
        cpu_3_data_master_read_last_time <= cpu_3_data_master_read;
    end


  //cpu_3_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_3_data_master_read != cpu_3_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_3_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_3_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_write_last_time <= 0;
      else 
        cpu_3_data_master_write_last_time <= cpu_3_data_master_write;
    end


  //cpu_3_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_3_data_master_write != cpu_3_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_3_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_3_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_writedata_last_time <= 0;
      else 
        cpu_3_data_master_writedata_last_time <= cpu_3_data_master_writedata;
    end


  //cpu_3_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_3_data_master_writedata != cpu_3_data_master_writedata_last_time) & cpu_3_data_master_write)
        begin
          $write("%0d ns: cpu_3_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_3_instruction_master_arbitrator (
                                             // inputs:
                                              clk,
                                              cpu_3_instruction_master_address,
                                              cpu_3_instruction_master_granted_cpu_3_jtag_debug_module,
                                              cpu_3_instruction_master_granted_nios_system_clock_6_in,
                                              cpu_3_instruction_master_granted_onchip_memory2_0_s1,
                                              cpu_3_instruction_master_granted_onchip_memory2_1_s1,
                                              cpu_3_instruction_master_granted_onchip_memory2_2_s1,
                                              cpu_3_instruction_master_granted_onchip_memory2_3_s1,
                                              cpu_3_instruction_master_granted_sram_0_avalon_sram_slave,
                                              cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module,
                                              cpu_3_instruction_master_qualified_request_nios_system_clock_6_in,
                                              cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1,
                                              cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1,
                                              cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1,
                                              cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1,
                                              cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave,
                                              cpu_3_instruction_master_read,
                                              cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module,
                                              cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in,
                                              cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1,
                                              cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1,
                                              cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1,
                                              cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1,
                                              cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave,
                                              cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                              cpu_3_instruction_master_requests_cpu_3_jtag_debug_module,
                                              cpu_3_instruction_master_requests_nios_system_clock_6_in,
                                              cpu_3_instruction_master_requests_onchip_memory2_0_s1,
                                              cpu_3_instruction_master_requests_onchip_memory2_1_s1,
                                              cpu_3_instruction_master_requests_onchip_memory2_2_s1,
                                              cpu_3_instruction_master_requests_onchip_memory2_3_s1,
                                              cpu_3_instruction_master_requests_sram_0_avalon_sram_slave,
                                              cpu_3_jtag_debug_module_readdata_from_sa,
                                              d1_cpu_3_jtag_debug_module_end_xfer,
                                              d1_nios_system_clock_6_in_end_xfer,
                                              d1_onchip_memory2_0_s1_end_xfer,
                                              d1_onchip_memory2_1_s1_end_xfer,
                                              d1_onchip_memory2_2_s1_end_xfer,
                                              d1_onchip_memory2_3_s1_end_xfer,
                                              d1_sram_0_avalon_sram_slave_end_xfer,
                                              nios_system_clock_6_in_readdata_from_sa,
                                              nios_system_clock_6_in_waitrequest_from_sa,
                                              onchip_memory2_0_s1_readdata_from_sa,
                                              onchip_memory2_1_s1_readdata_from_sa,
                                              onchip_memory2_2_s1_readdata_from_sa,
                                              onchip_memory2_3_s1_readdata_from_sa,
                                              reset_n,
                                              sram_0_avalon_sram_slave_readdata_from_sa,

                                             // outputs:
                                              cpu_3_instruction_master_address_to_slave,
                                              cpu_3_instruction_master_dbs_address,
                                              cpu_3_instruction_master_latency_counter,
                                              cpu_3_instruction_master_readdata,
                                              cpu_3_instruction_master_readdatavalid,
                                              cpu_3_instruction_master_waitrequest
                                           )
;

  output  [ 24: 0] cpu_3_instruction_master_address_to_slave;
  output  [  1: 0] cpu_3_instruction_master_dbs_address;
  output           cpu_3_instruction_master_latency_counter;
  output  [ 31: 0] cpu_3_instruction_master_readdata;
  output           cpu_3_instruction_master_readdatavalid;
  output           cpu_3_instruction_master_waitrequest;
  input            clk;
  input   [ 24: 0] cpu_3_instruction_master_address;
  input            cpu_3_instruction_master_granted_cpu_3_jtag_debug_module;
  input            cpu_3_instruction_master_granted_nios_system_clock_6_in;
  input            cpu_3_instruction_master_granted_onchip_memory2_0_s1;
  input            cpu_3_instruction_master_granted_onchip_memory2_1_s1;
  input            cpu_3_instruction_master_granted_onchip_memory2_2_s1;
  input            cpu_3_instruction_master_granted_onchip_memory2_3_s1;
  input            cpu_3_instruction_master_granted_sram_0_avalon_sram_slave;
  input            cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module;
  input            cpu_3_instruction_master_qualified_request_nios_system_clock_6_in;
  input            cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1;
  input            cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1;
  input            cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1;
  input            cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1;
  input            cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  input            cpu_3_instruction_master_read;
  input            cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module;
  input            cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in;
  input            cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1;
  input            cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1;
  input            cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1;
  input            cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1;
  input            cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  input            cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_instruction_master_requests_cpu_3_jtag_debug_module;
  input            cpu_3_instruction_master_requests_nios_system_clock_6_in;
  input            cpu_3_instruction_master_requests_onchip_memory2_0_s1;
  input            cpu_3_instruction_master_requests_onchip_memory2_1_s1;
  input            cpu_3_instruction_master_requests_onchip_memory2_2_s1;
  input            cpu_3_instruction_master_requests_onchip_memory2_3_s1;
  input            cpu_3_instruction_master_requests_sram_0_avalon_sram_slave;
  input   [ 31: 0] cpu_3_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_3_jtag_debug_module_end_xfer;
  input            d1_nios_system_clock_6_in_end_xfer;
  input            d1_onchip_memory2_0_s1_end_xfer;
  input            d1_onchip_memory2_1_s1_end_xfer;
  input            d1_onchip_memory2_2_s1_end_xfer;
  input            d1_onchip_memory2_3_s1_end_xfer;
  input            d1_sram_0_avalon_sram_slave_end_xfer;
  input   [ 15: 0] nios_system_clock_6_in_readdata_from_sa;
  input            nios_system_clock_6_in_waitrequest_from_sa;
  input   [ 31: 0] onchip_memory2_0_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_1_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_2_s1_readdata_from_sa;
  input   [ 31: 0] onchip_memory2_3_s1_readdata_from_sa;
  input            reset_n;
  input   [ 15: 0] sram_0_avalon_sram_slave_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] cpu_3_instruction_master_address_last_time;
  wire    [ 24: 0] cpu_3_instruction_master_address_to_slave;
  reg     [  1: 0] cpu_3_instruction_master_dbs_address;
  wire    [  1: 0] cpu_3_instruction_master_dbs_increment;
  reg     [  1: 0] cpu_3_instruction_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_3_instruction_master_dbs_rdv_counter_inc;
  wire             cpu_3_instruction_master_is_granted_some_slave;
  reg              cpu_3_instruction_master_latency_counter;
  wire    [  1: 0] cpu_3_instruction_master_next_dbs_rdv_counter;
  reg              cpu_3_instruction_master_read_but_no_slave_selected;
  reg              cpu_3_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_3_instruction_master_readdata;
  wire             cpu_3_instruction_master_readdatavalid;
  wire             cpu_3_instruction_master_run;
  wire             cpu_3_instruction_master_waitrequest;
  reg     [ 15: 0] dbs_16_reg_segment_0;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire             p1_cpu_3_instruction_master_latency_counter;
  wire    [ 15: 0] p1_dbs_16_reg_segment_0;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_3_instruction_master_readdatavalid;
  wire             r_0;
  wire             r_2;
  wire             r_3;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module | ~cpu_3_instruction_master_requests_cpu_3_jtag_debug_module) & (cpu_3_instruction_master_granted_cpu_3_jtag_debug_module | ~cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module) & ((~cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module | ~cpu_3_instruction_master_read | (1 & ~d1_cpu_3_jtag_debug_module_end_xfer & cpu_3_instruction_master_read)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_3_instruction_master_run = r_0 & r_2 & r_3;

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_3_instruction_master_qualified_request_nios_system_clock_6_in | ~cpu_3_instruction_master_requests_nios_system_clock_6_in) & ((~cpu_3_instruction_master_qualified_request_nios_system_clock_6_in | ~cpu_3_instruction_master_read | (1 & ~nios_system_clock_6_in_waitrequest_from_sa & (cpu_3_instruction_master_dbs_address[1]) & cpu_3_instruction_master_read))) & 1 & (cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1 | ~cpu_3_instruction_master_requests_onchip_memory2_0_s1) & (cpu_3_instruction_master_granted_onchip_memory2_0_s1 | ~cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1) & ((~cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1 | ~(cpu_3_instruction_master_read) | (1 & (cpu_3_instruction_master_read)))) & 1 & (cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1 | ~cpu_3_instruction_master_requests_onchip_memory2_1_s1) & (cpu_3_instruction_master_granted_onchip_memory2_1_s1 | ~cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1) & ((~cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1 | ~(cpu_3_instruction_master_read) | (1 & (cpu_3_instruction_master_read)))) & 1 & (cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1 | ~cpu_3_instruction_master_requests_onchip_memory2_2_s1) & (cpu_3_instruction_master_granted_onchip_memory2_2_s1 | ~cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1) & ((~cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1 | ~(cpu_3_instruction_master_read) | (1 & (cpu_3_instruction_master_read))));

  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1 | ~cpu_3_instruction_master_requests_onchip_memory2_3_s1) & (cpu_3_instruction_master_granted_onchip_memory2_3_s1 | ~cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1) & ((~cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1 | ~(cpu_3_instruction_master_read) | (1 & (cpu_3_instruction_master_read)))) & 1 & (cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_3_instruction_master_requests_sram_0_avalon_sram_slave) & (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave | ~cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave) & ((~cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave | ~cpu_3_instruction_master_read | (1 & (cpu_3_instruction_master_dbs_address[1]) & cpu_3_instruction_master_read)));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_3_instruction_master_address_to_slave = cpu_3_instruction_master_address[24 : 0];

  //cpu_3_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_3_instruction_master_read_but_no_slave_selected <= cpu_3_instruction_master_read & cpu_3_instruction_master_run & ~cpu_3_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_3_instruction_master_is_granted_some_slave = cpu_3_instruction_master_granted_cpu_3_jtag_debug_module |
    cpu_3_instruction_master_granted_nios_system_clock_6_in |
    cpu_3_instruction_master_granted_onchip_memory2_0_s1 |
    cpu_3_instruction_master_granted_onchip_memory2_1_s1 |
    cpu_3_instruction_master_granted_onchip_memory2_2_s1 |
    cpu_3_instruction_master_granted_onchip_memory2_3_s1 |
    cpu_3_instruction_master_granted_sram_0_avalon_sram_slave;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_3_instruction_master_readdatavalid = cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1 |
    cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1 |
    cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1 |
    cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1 |
    (cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave & dbs_rdv_counter_overflow);

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_3_instruction_master_readdatavalid = cpu_3_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_3_instruction_master_readdatavalid |
    cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module |
    cpu_3_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_3_instruction_master_readdatavalid |
    (cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in & dbs_counter_overflow) |
    cpu_3_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_3_instruction_master_readdatavalid |
    cpu_3_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_3_instruction_master_readdatavalid |
    cpu_3_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_3_instruction_master_readdatavalid |
    cpu_3_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_3_instruction_master_readdatavalid |
    cpu_3_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_3_instruction_master_readdatavalid;

  //cpu_3/instruction_master readdata mux, which is an e_mux
  assign cpu_3_instruction_master_readdata = ({32 {~(cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module & cpu_3_instruction_master_read)}} | cpu_3_jtag_debug_module_readdata_from_sa) &
    ({32 {~(cpu_3_instruction_master_qualified_request_nios_system_clock_6_in & cpu_3_instruction_master_read)}} | {nios_system_clock_6_in_readdata_from_sa[15 : 0],
    dbs_16_reg_segment_0}) &
    ({32 {~cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1}} | onchip_memory2_0_s1_readdata_from_sa) &
    ({32 {~cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1}} | onchip_memory2_1_s1_readdata_from_sa) &
    ({32 {~cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1}} | onchip_memory2_2_s1_readdata_from_sa) &
    ({32 {~cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1}} | onchip_memory2_3_s1_readdata_from_sa) &
    ({32 {~cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave}} | {sram_0_avalon_sram_slave_readdata_from_sa[15 : 0],
    dbs_latent_16_reg_segment_0});

  //actual waitrequest port, which is an e_assign
  assign cpu_3_instruction_master_waitrequest = ~cpu_3_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_instruction_master_latency_counter <= 0;
      else 
        cpu_3_instruction_master_latency_counter <= p1_cpu_3_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_3_instruction_master_latency_counter = ((cpu_3_instruction_master_run & cpu_3_instruction_master_read))? latency_load_value :
    (cpu_3_instruction_master_latency_counter)? cpu_3_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = ({1 {cpu_3_instruction_master_requests_onchip_memory2_0_s1}} & 1) |
    ({1 {cpu_3_instruction_master_requests_onchip_memory2_1_s1}} & 1) |
    ({1 {cpu_3_instruction_master_requests_onchip_memory2_2_s1}} & 1) |
    ({1 {cpu_3_instruction_master_requests_onchip_memory2_3_s1}} & 1);

  //input to dbs-16 stored 0, which is an e_mux
  assign p1_dbs_16_reg_segment_0 = nios_system_clock_6_in_readdata_from_sa;

  //dbs register for dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_16_reg_segment_0 <= 0;
      else if (dbs_count_enable & ((cpu_3_instruction_master_dbs_address[1]) == 0))
          dbs_16_reg_segment_0 <= p1_dbs_16_reg_segment_0;
    end


  //dbs count increment, which is an e_mux
  assign cpu_3_instruction_master_dbs_increment = (cpu_3_instruction_master_requests_nios_system_clock_6_in)? 2 :
    (cpu_3_instruction_master_requests_sram_0_avalon_sram_slave)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_3_instruction_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_3_instruction_master_dbs_address + cpu_3_instruction_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_instruction_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_3_instruction_master_dbs_address <= next_dbs_address;
    end


  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (cpu_3_instruction_master_granted_nios_system_clock_6_in & cpu_3_instruction_master_read & 1 & 1 & ~nios_system_clock_6_in_waitrequest_from_sa) |
    (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave & cpu_3_instruction_master_read & 1 & 1);

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = sram_0_avalon_sram_slave_readdata_from_sa;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_3_instruction_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_3_instruction_master_next_dbs_rdv_counter = cpu_3_instruction_master_dbs_rdv_counter + cpu_3_instruction_master_dbs_rdv_counter_inc;

  //cpu_3_instruction_master_rdv_inc_mux, which is an e_mux
  assign cpu_3_instruction_master_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_instruction_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_3_instruction_master_dbs_rdv_counter <= cpu_3_instruction_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_3_instruction_master_dbs_rdv_counter[1] & ~cpu_3_instruction_master_next_dbs_rdv_counter[1];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_3_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_instruction_master_address_last_time <= 0;
      else 
        cpu_3_instruction_master_address_last_time <= cpu_3_instruction_master_address;
    end


  //cpu_3/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_3_instruction_master_waitrequest & (cpu_3_instruction_master_read);
    end


  //cpu_3_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_3_instruction_master_address != cpu_3_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_3_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_3_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_instruction_master_read_last_time <= 0;
      else 
        cpu_3_instruction_master_read_last_time <= cpu_3_instruction_master_read;
    end


  //cpu_3_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_3_instruction_master_read != cpu_3_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_3_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_3_altera_nios_custom_instr_floating_point_inst_s1_arbitrator (
                                                                          // inputs:
                                                                           clk,
                                                                           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done,
                                                                           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result,
                                                                           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select,
                                                                           cpu_3_custom_instruction_master_multi_clk_en,
                                                                           cpu_3_custom_instruction_master_multi_dataa,
                                                                           cpu_3_custom_instruction_master_multi_datab,
                                                                           cpu_3_custom_instruction_master_multi_n,
                                                                           cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1,
                                                                           reset_n,

                                                                          // outputs:
                                                                           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_clk_en,
                                                                           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_dataa,
                                                                           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_datab,
                                                                           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa,
                                                                           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_n,
                                                                           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_reset,
                                                                           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa,
                                                                           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_start
                                                                        )
;

  output           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  output  [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  output  [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_datab;
  output           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  output  [  1: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_n;
  output           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_reset;
  output  [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  output           cpu_3_altera_nios_custom_instr_floating_point_inst_s1_start;
  input            clk;
  input            cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done;
  input   [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result;
  input            cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select;
  input            cpu_3_custom_instruction_master_multi_clk_en;
  input   [ 31: 0] cpu_3_custom_instruction_master_multi_dataa;
  input   [ 31: 0] cpu_3_custom_instruction_master_multi_datab;
  input   [  7: 0] cpu_3_custom_instruction_master_multi_n;
  input            cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1;
  input            reset_n;

  wire             cpu_3_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  wire    [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  wire    [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_datab;
  wire             cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  wire    [  1: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_n;
  wire             cpu_3_altera_nios_custom_instr_floating_point_inst_s1_reset;
  wire    [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  wire             cpu_3_altera_nios_custom_instr_floating_point_inst_s1_start;
  assign cpu_3_altera_nios_custom_instr_floating_point_inst_s1_clk_en = cpu_3_custom_instruction_master_multi_clk_en;
  assign cpu_3_altera_nios_custom_instr_floating_point_inst_s1_dataa = cpu_3_custom_instruction_master_multi_dataa;
  assign cpu_3_altera_nios_custom_instr_floating_point_inst_s1_datab = cpu_3_custom_instruction_master_multi_datab;
  assign cpu_3_altera_nios_custom_instr_floating_point_inst_s1_n = cpu_3_custom_instruction_master_multi_n;
  assign cpu_3_altera_nios_custom_instr_floating_point_inst_s1_start = cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1;
  //assign cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa = cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa = cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result;

  //assign cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa = cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa = cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done;

  //cpu_3_altera_nios_custom_instr_floating_point_inst/s1 local reset_n, which is an e_assign
  assign cpu_3_altera_nios_custom_instr_floating_point_inst_s1_reset = ~reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_0_avalon_jtag_slave_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   cpu_0_data_master_address_to_slave,
                                                   cpu_0_data_master_latency_counter,
                                                   cpu_0_data_master_read,
                                                   cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                   cpu_0_data_master_write,
                                                   cpu_0_data_master_writedata,
                                                   jtag_uart_0_avalon_jtag_slave_dataavailable,
                                                   jtag_uart_0_avalon_jtag_slave_irq,
                                                   jtag_uart_0_avalon_jtag_slave_readdata,
                                                   jtag_uart_0_avalon_jtag_slave_readyfordata,
                                                   jtag_uart_0_avalon_jtag_slave_waitrequest,
                                                   reset_n,

                                                  // outputs:
                                                   cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave,
                                                   cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave,
                                                   cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave,
                                                   cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave,
                                                   d1_jtag_uart_0_avalon_jtag_slave_end_xfer,
                                                   jtag_uart_0_avalon_jtag_slave_address,
                                                   jtag_uart_0_avalon_jtag_slave_chipselect,
                                                   jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_irq_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_read_n,
                                                   jtag_uart_0_avalon_jtag_slave_readdata_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_reset_n,
                                                   jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_write_n,
                                                   jtag_uart_0_avalon_jtag_slave_writedata
                                                )
;

  output           cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave;
  output           cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave;
  output           cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  output           cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;
  output           d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  output           jtag_uart_0_avalon_jtag_slave_address;
  output           jtag_uart_0_avalon_jtag_slave_chipselect;
  output           jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_reset_n;
  output           jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_0_avalon_jtag_slave_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input            jtag_uart_0_avalon_jtag_slave_dataavailable;
  input            jtag_uart_0_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata;
  input            jtag_uart_0_avalon_jtag_slave_readyfordata;
  input            jtag_uart_0_avalon_jtag_slave_waitrequest;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_saved_grant_jtag_uart_0_avalon_jtag_slave;
  reg              d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_address;
  wire             jtag_uart_0_avalon_jtag_slave_allgrants;
  wire             jtag_uart_0_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_0_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_0_avalon_jtag_slave_arb_counter_enable;
  reg     [  2: 0] jtag_uart_0_avalon_jtag_slave_arb_share_counter;
  wire    [  2: 0] jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
  wire    [  2: 0] jtag_uart_0_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_0_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_0_avalon_jtag_slave_chipselect;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_0_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_0_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_0_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_0_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_0_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_0_avalon_jtag_slave_reset_n;
  reg              jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_0_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_0_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_writedata;
  wire    [ 24: 0] shifted_address_to_jtag_uart_0_avalon_jtag_slave_from_cpu_0_data_master;
  wire             wait_for_jtag_uart_0_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_0_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_0_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave));
  //assign jtag_uart_0_avalon_jtag_slave_readdata_from_sa = jtag_uart_0_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_readdata_from_sa = jtag_uart_0_avalon_jtag_slave_readdata;

  assign cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave = ({cpu_0_data_master_address_to_slave[24 : 3] , 3'b0} == 25'h19030c8) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //assign jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_0_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_0_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_0_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_0_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_0_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_0_avalon_jtag_slave_waitrequest;

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_arb_share_set_values = 1;

  //jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests = cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;

  //jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant = 0;

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_0_avalon_jtag_slave_firsttransfer ? (jtag_uart_0_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_0_avalon_jtag_slave_arb_share_counter ? (jtag_uart_0_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_0_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_allgrants = |jtag_uart_0_avalon_jtag_slave_grant_vector;

  //jtag_uart_0_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_end_xfer = ~(jtag_uart_0_avalon_jtag_slave_waits_for_read | jtag_uart_0_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave = jtag_uart_0_avalon_jtag_slave_end_xfer & (~jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave & jtag_uart_0_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave & ~jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_0_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_0_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_0_avalon_jtag_slave_arb_share_counter <= jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_0_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave & ~jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //cpu_0/data_master jtag_uart_0/avalon_jtag_slave arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;

  //cpu_0/data_master jtag_uart_0/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //jtag_uart_0_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_any_continuerequest = 1;

  //cpu_0_data_master_continuerequest continued request, which is an e_assign
  assign cpu_0_data_master_continuerequest = 1;

  assign cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave = cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))));
  //local readdatavalid cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave, which is an e_mux
  assign cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave = cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_read & ~jtag_uart_0_avalon_jtag_slave_waits_for_read;

  //jtag_uart_0_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_writedata = cpu_0_data_master_writedata;

  //master is always granted when requested
  assign cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave = cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave;

  //cpu_0/data_master saved-grant jtag_uart_0/avalon_jtag_slave, which is an e_assign
  assign cpu_0_data_master_saved_grant_jtag_uart_0_avalon_jtag_slave = cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart_0/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_0_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_0_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_0_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_0_avalon_jtag_slave_chipselect = cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave;
  //jtag_uart_0_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_firsttransfer = jtag_uart_0_avalon_jtag_slave_begins_xfer ? jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_0_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_0_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_0_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_0_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_0_avalon_jtag_slave_begins_xfer)
          jtag_uart_0_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_0_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_0_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_read_n = ~(cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_read);

  //~jtag_uart_0_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_write_n = ~(cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_write);

  assign shifted_address_to_jtag_uart_0_avalon_jtag_slave_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //jtag_uart_0_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_address = shifted_address_to_jtag_uart_0_avalon_jtag_slave_from_cpu_0_data_master >> 2;

  //d1_jtag_uart_0_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_0_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_0_avalon_jtag_slave_end_xfer <= jtag_uart_0_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_0_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_waits_for_read = jtag_uart_0_avalon_jtag_slave_in_a_read_cycle & jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_0_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_in_a_read_cycle = cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_0_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_0_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_waits_for_write = jtag_uart_0_avalon_jtag_slave_in_a_write_cycle & jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_0_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_in_a_write_cycle = cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_0_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_0_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_0_avalon_jtag_slave_irq_from_sa = jtag_uart_0_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_irq_from_sa = jtag_uart_0_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart_0/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_1_avalon_jtag_slave_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   cpu_1_data_master_address_to_slave,
                                                   cpu_1_data_master_latency_counter,
                                                   cpu_1_data_master_read,
                                                   cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                   cpu_1_data_master_write,
                                                   cpu_1_data_master_writedata,
                                                   jtag_uart_1_avalon_jtag_slave_dataavailable,
                                                   jtag_uart_1_avalon_jtag_slave_irq,
                                                   jtag_uart_1_avalon_jtag_slave_readdata,
                                                   jtag_uart_1_avalon_jtag_slave_readyfordata,
                                                   jtag_uart_1_avalon_jtag_slave_waitrequest,
                                                   reset_n,

                                                  // outputs:
                                                   cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave,
                                                   cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave,
                                                   cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave,
                                                   cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave,
                                                   d1_jtag_uart_1_avalon_jtag_slave_end_xfer,
                                                   jtag_uart_1_avalon_jtag_slave_address,
                                                   jtag_uart_1_avalon_jtag_slave_chipselect,
                                                   jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa,
                                                   jtag_uart_1_avalon_jtag_slave_irq_from_sa,
                                                   jtag_uart_1_avalon_jtag_slave_read_n,
                                                   jtag_uart_1_avalon_jtag_slave_readdata_from_sa,
                                                   jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa,
                                                   jtag_uart_1_avalon_jtag_slave_reset_n,
                                                   jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa,
                                                   jtag_uart_1_avalon_jtag_slave_write_n,
                                                   jtag_uart_1_avalon_jtag_slave_writedata
                                                )
;

  output           cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave;
  output           cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave;
  output           cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave;
  output           cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave;
  output           d1_jtag_uart_1_avalon_jtag_slave_end_xfer;
  output           jtag_uart_1_avalon_jtag_slave_address;
  output           jtag_uart_1_avalon_jtag_slave_chipselect;
  output           jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_1_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_1_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_1_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_1_avalon_jtag_slave_reset_n;
  output           jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_1_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_1_avalon_jtag_slave_writedata;
  input            clk;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input            jtag_uart_1_avalon_jtag_slave_dataavailable;
  input            jtag_uart_1_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_1_avalon_jtag_slave_readdata;
  input            jtag_uart_1_avalon_jtag_slave_readyfordata;
  input            jtag_uart_1_avalon_jtag_slave_waitrequest;
  input            reset_n;

  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave;
  wire             cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave;
  wire             cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave;
  wire             cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave;
  wire             cpu_1_data_master_saved_grant_jtag_uart_1_avalon_jtag_slave;
  reg              d1_jtag_uart_1_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_1_avalon_jtag_slave_address;
  wire             jtag_uart_1_avalon_jtag_slave_allgrants;
  wire             jtag_uart_1_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_1_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_1_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_1_avalon_jtag_slave_arb_counter_enable;
  reg     [  2: 0] jtag_uart_1_avalon_jtag_slave_arb_share_counter;
  wire    [  2: 0] jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value;
  wire    [  2: 0] jtag_uart_1_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_1_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_1_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_1_avalon_jtag_slave_chipselect;
  wire             jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_1_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_1_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_1_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_1_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_1_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_1_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_1_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_1_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_1_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_1_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_1_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_1_avalon_jtag_slave_reset_n;
  reg              jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_1_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_1_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_1_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_1_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_1_avalon_jtag_slave_writedata;
  wire    [ 24: 0] shifted_address_to_jtag_uart_1_avalon_jtag_slave_from_cpu_1_data_master;
  wire             wait_for_jtag_uart_1_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_1_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_1_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave));
  //assign jtag_uart_1_avalon_jtag_slave_readdata_from_sa = jtag_uart_1_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_readdata_from_sa = jtag_uart_1_avalon_jtag_slave_readdata;

  assign cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave = ({cpu_1_data_master_address_to_slave[24 : 3] , 3'b0} == 25'h60) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //assign jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_1_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_1_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_1_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_1_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_1_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_1_avalon_jtag_slave_waitrequest;

  //jtag_uart_1_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_1_avalon_jtag_slave_arb_share_set_values = 1;

  //jtag_uart_1_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_1_avalon_jtag_slave_non_bursting_master_requests = cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave;

  //jtag_uart_1_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_1_avalon_jtag_slave_any_bursting_master_saved_grant = 0;

  //jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_1_avalon_jtag_slave_firsttransfer ? (jtag_uart_1_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_1_avalon_jtag_slave_arb_share_counter ? (jtag_uart_1_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_1_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_1_avalon_jtag_slave_allgrants = |jtag_uart_1_avalon_jtag_slave_grant_vector;

  //jtag_uart_1_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_end_xfer = ~(jtag_uart_1_avalon_jtag_slave_waits_for_read | jtag_uart_1_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave = jtag_uart_1_avalon_jtag_slave_end_xfer & (~jtag_uart_1_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_1_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave & jtag_uart_1_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave & ~jtag_uart_1_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_1_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_1_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_1_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_1_avalon_jtag_slave_arb_share_counter <= jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_1_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_1_avalon_jtag_slave & ~jtag_uart_1_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //cpu_1/data_master jtag_uart_1/avalon_jtag_slave arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_1_avalon_jtag_slave_arb_share_counter_next_value;

  //cpu_1/data_master jtag_uart_1/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //jtag_uart_1_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_any_continuerequest = 1;

  //cpu_1_data_master_continuerequest continued request, which is an e_assign
  assign cpu_1_data_master_continuerequest = 1;

  assign cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave = cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave & ~((cpu_1_data_master_read & ((cpu_1_data_master_latency_counter != 0) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))));
  //local readdatavalid cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave, which is an e_mux
  assign cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave = cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave & cpu_1_data_master_read & ~jtag_uart_1_avalon_jtag_slave_waits_for_read;

  //jtag_uart_1_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_1_avalon_jtag_slave_writedata = cpu_1_data_master_writedata;

  //master is always granted when requested
  assign cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave = cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave;

  //cpu_1/data_master saved-grant jtag_uart_1/avalon_jtag_slave, which is an e_assign
  assign cpu_1_data_master_saved_grant_jtag_uart_1_avalon_jtag_slave = cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart_1/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_1_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_1_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_1_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_1_avalon_jtag_slave_chipselect = cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave;
  //jtag_uart_1_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_firsttransfer = jtag_uart_1_avalon_jtag_slave_begins_xfer ? jtag_uart_1_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_1_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_1_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_1_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_1_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_1_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_1_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_1_avalon_jtag_slave_begins_xfer)
          jtag_uart_1_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_1_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_1_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_1_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_1_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_1_avalon_jtag_slave_read_n = ~(cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave & cpu_1_data_master_read);

  //~jtag_uart_1_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_1_avalon_jtag_slave_write_n = ~(cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave & cpu_1_data_master_write);

  assign shifted_address_to_jtag_uart_1_avalon_jtag_slave_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  //jtag_uart_1_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_1_avalon_jtag_slave_address = shifted_address_to_jtag_uart_1_avalon_jtag_slave_from_cpu_1_data_master >> 2;

  //d1_jtag_uart_1_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_1_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_1_avalon_jtag_slave_end_xfer <= jtag_uart_1_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_1_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_1_avalon_jtag_slave_waits_for_read = jtag_uart_1_avalon_jtag_slave_in_a_read_cycle & jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_1_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_in_a_read_cycle = cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave & cpu_1_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_1_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_1_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_1_avalon_jtag_slave_waits_for_write = jtag_uart_1_avalon_jtag_slave_in_a_write_cycle & jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_1_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_in_a_write_cycle = cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave & cpu_1_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_1_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_1_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_1_avalon_jtag_slave_irq_from_sa = jtag_uart_1_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_1_avalon_jtag_slave_irq_from_sa = jtag_uart_1_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart_1/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_2_avalon_jtag_slave_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   cpu_2_data_master_address_to_slave,
                                                   cpu_2_data_master_latency_counter,
                                                   cpu_2_data_master_read,
                                                   cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                   cpu_2_data_master_write,
                                                   cpu_2_data_master_writedata,
                                                   jtag_uart_2_avalon_jtag_slave_dataavailable,
                                                   jtag_uart_2_avalon_jtag_slave_irq,
                                                   jtag_uart_2_avalon_jtag_slave_readdata,
                                                   jtag_uart_2_avalon_jtag_slave_readyfordata,
                                                   jtag_uart_2_avalon_jtag_slave_waitrequest,
                                                   reset_n,

                                                  // outputs:
                                                   cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave,
                                                   cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave,
                                                   cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave,
                                                   cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave,
                                                   d1_jtag_uart_2_avalon_jtag_slave_end_xfer,
                                                   jtag_uart_2_avalon_jtag_slave_address,
                                                   jtag_uart_2_avalon_jtag_slave_chipselect,
                                                   jtag_uart_2_avalon_jtag_slave_dataavailable_from_sa,
                                                   jtag_uart_2_avalon_jtag_slave_irq_from_sa,
                                                   jtag_uart_2_avalon_jtag_slave_read_n,
                                                   jtag_uart_2_avalon_jtag_slave_readdata_from_sa,
                                                   jtag_uart_2_avalon_jtag_slave_readyfordata_from_sa,
                                                   jtag_uart_2_avalon_jtag_slave_reset_n,
                                                   jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa,
                                                   jtag_uart_2_avalon_jtag_slave_write_n,
                                                   jtag_uart_2_avalon_jtag_slave_writedata
                                                )
;

  output           cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave;
  output           cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave;
  output           cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave;
  output           cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave;
  output           d1_jtag_uart_2_avalon_jtag_slave_end_xfer;
  output           jtag_uart_2_avalon_jtag_slave_address;
  output           jtag_uart_2_avalon_jtag_slave_chipselect;
  output           jtag_uart_2_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_2_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_2_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_2_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_2_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_2_avalon_jtag_slave_reset_n;
  output           jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_2_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_2_avalon_jtag_slave_writedata;
  input            clk;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input            jtag_uart_2_avalon_jtag_slave_dataavailable;
  input            jtag_uart_2_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_2_avalon_jtag_slave_readdata;
  input            jtag_uart_2_avalon_jtag_slave_readyfordata;
  input            jtag_uart_2_avalon_jtag_slave_waitrequest;
  input            reset_n;

  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave;
  wire             cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave;
  wire             cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave;
  wire             cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave;
  wire             cpu_2_data_master_saved_grant_jtag_uart_2_avalon_jtag_slave;
  reg              d1_jtag_uart_2_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_2_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_2_avalon_jtag_slave_address;
  wire             jtag_uart_2_avalon_jtag_slave_allgrants;
  wire             jtag_uart_2_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_2_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_2_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_2_avalon_jtag_slave_arb_counter_enable;
  reg     [  2: 0] jtag_uart_2_avalon_jtag_slave_arb_share_counter;
  wire    [  2: 0] jtag_uart_2_avalon_jtag_slave_arb_share_counter_next_value;
  wire    [  2: 0] jtag_uart_2_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_2_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_2_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_2_avalon_jtag_slave_chipselect;
  wire             jtag_uart_2_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_2_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_2_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_2_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_2_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_2_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_2_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_2_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_2_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_2_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_2_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_2_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_2_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_2_avalon_jtag_slave_reset_n;
  reg              jtag_uart_2_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_2_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_2_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_2_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_2_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_2_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_2_avalon_jtag_slave_writedata;
  wire    [ 24: 0] shifted_address_to_jtag_uart_2_avalon_jtag_slave_from_cpu_2_data_master;
  wire             wait_for_jtag_uart_2_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_2_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_2_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave));
  //assign jtag_uart_2_avalon_jtag_slave_readdata_from_sa = jtag_uart_2_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_readdata_from_sa = jtag_uart_2_avalon_jtag_slave_readdata;

  assign cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave = ({cpu_2_data_master_address_to_slave[24 : 3] , 3'b0} == 25'h68) & (cpu_2_data_master_read | cpu_2_data_master_write);
  //assign jtag_uart_2_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_2_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_2_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_2_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_2_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_2_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_2_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_2_avalon_jtag_slave_waitrequest;

  //jtag_uart_2_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_2_avalon_jtag_slave_arb_share_set_values = 1;

  //jtag_uart_2_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_2_avalon_jtag_slave_non_bursting_master_requests = cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave;

  //jtag_uart_2_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_2_avalon_jtag_slave_any_bursting_master_saved_grant = 0;

  //jtag_uart_2_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_2_avalon_jtag_slave_firsttransfer ? (jtag_uart_2_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_2_avalon_jtag_slave_arb_share_counter ? (jtag_uart_2_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_2_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_2_avalon_jtag_slave_allgrants = |jtag_uart_2_avalon_jtag_slave_grant_vector;

  //jtag_uart_2_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_end_xfer = ~(jtag_uart_2_avalon_jtag_slave_waits_for_read | jtag_uart_2_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_2_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_2_avalon_jtag_slave = jtag_uart_2_avalon_jtag_slave_end_xfer & (~jtag_uart_2_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_2_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_2_avalon_jtag_slave & jtag_uart_2_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_2_avalon_jtag_slave & ~jtag_uart_2_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_2_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_2_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_2_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_2_avalon_jtag_slave_arb_share_counter <= jtag_uart_2_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_2_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_2_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_2_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_2_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_2_avalon_jtag_slave & ~jtag_uart_2_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_2_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_2_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //cpu_2/data_master jtag_uart_2/avalon_jtag_slave arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = jtag_uart_2_avalon_jtag_slave_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //jtag_uart_2_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_2_avalon_jtag_slave_arb_share_counter_next_value;

  //cpu_2/data_master jtag_uart_2/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = jtag_uart_2_avalon_jtag_slave_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //jtag_uart_2_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_any_continuerequest = 1;

  //cpu_2_data_master_continuerequest continued request, which is an e_assign
  assign cpu_2_data_master_continuerequest = 1;

  assign cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave = cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave & ~((cpu_2_data_master_read & ((cpu_2_data_master_latency_counter != 0) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))));
  //local readdatavalid cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave, which is an e_mux
  assign cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave = cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave & cpu_2_data_master_read & ~jtag_uart_2_avalon_jtag_slave_waits_for_read;

  //jtag_uart_2_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_2_avalon_jtag_slave_writedata = cpu_2_data_master_writedata;

  //master is always granted when requested
  assign cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave = cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave;

  //cpu_2/data_master saved-grant jtag_uart_2/avalon_jtag_slave, which is an e_assign
  assign cpu_2_data_master_saved_grant_jtag_uart_2_avalon_jtag_slave = cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart_2/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_2_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_2_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_2_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_2_avalon_jtag_slave_chipselect = cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave;
  //jtag_uart_2_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_firsttransfer = jtag_uart_2_avalon_jtag_slave_begins_xfer ? jtag_uart_2_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_2_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_2_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_2_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_2_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_2_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_2_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_2_avalon_jtag_slave_begins_xfer)
          jtag_uart_2_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_2_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_2_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_2_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_2_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_2_avalon_jtag_slave_read_n = ~(cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave & cpu_2_data_master_read);

  //~jtag_uart_2_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_2_avalon_jtag_slave_write_n = ~(cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave & cpu_2_data_master_write);

  assign shifted_address_to_jtag_uart_2_avalon_jtag_slave_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  //jtag_uart_2_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_2_avalon_jtag_slave_address = shifted_address_to_jtag_uart_2_avalon_jtag_slave_from_cpu_2_data_master >> 2;

  //d1_jtag_uart_2_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_2_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_2_avalon_jtag_slave_end_xfer <= jtag_uart_2_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_2_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_2_avalon_jtag_slave_waits_for_read = jtag_uart_2_avalon_jtag_slave_in_a_read_cycle & jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_2_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_in_a_read_cycle = cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave & cpu_2_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_2_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_2_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_2_avalon_jtag_slave_waits_for_write = jtag_uart_2_avalon_jtag_slave_in_a_write_cycle & jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_2_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_in_a_write_cycle = cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave & cpu_2_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_2_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_2_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_2_avalon_jtag_slave_irq_from_sa = jtag_uart_2_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_2_avalon_jtag_slave_irq_from_sa = jtag_uart_2_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart_2/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_3_avalon_jtag_slave_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   cpu_3_data_master_address_to_slave,
                                                   cpu_3_data_master_latency_counter,
                                                   cpu_3_data_master_read,
                                                   cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                   cpu_3_data_master_write,
                                                   cpu_3_data_master_writedata,
                                                   jtag_uart_3_avalon_jtag_slave_dataavailable,
                                                   jtag_uart_3_avalon_jtag_slave_irq,
                                                   jtag_uart_3_avalon_jtag_slave_readdata,
                                                   jtag_uart_3_avalon_jtag_slave_readyfordata,
                                                   jtag_uart_3_avalon_jtag_slave_waitrequest,
                                                   reset_n,

                                                  // outputs:
                                                   cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave,
                                                   cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave,
                                                   cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave,
                                                   cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave,
                                                   d1_jtag_uart_3_avalon_jtag_slave_end_xfer,
                                                   jtag_uart_3_avalon_jtag_slave_address,
                                                   jtag_uart_3_avalon_jtag_slave_chipselect,
                                                   jtag_uart_3_avalon_jtag_slave_dataavailable_from_sa,
                                                   jtag_uart_3_avalon_jtag_slave_irq_from_sa,
                                                   jtag_uart_3_avalon_jtag_slave_read_n,
                                                   jtag_uart_3_avalon_jtag_slave_readdata_from_sa,
                                                   jtag_uart_3_avalon_jtag_slave_readyfordata_from_sa,
                                                   jtag_uart_3_avalon_jtag_slave_reset_n,
                                                   jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa,
                                                   jtag_uart_3_avalon_jtag_slave_write_n,
                                                   jtag_uart_3_avalon_jtag_slave_writedata
                                                )
;

  output           cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave;
  output           cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave;
  output           cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave;
  output           cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave;
  output           d1_jtag_uart_3_avalon_jtag_slave_end_xfer;
  output           jtag_uart_3_avalon_jtag_slave_address;
  output           jtag_uart_3_avalon_jtag_slave_chipselect;
  output           jtag_uart_3_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_3_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_3_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_3_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_3_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_3_avalon_jtag_slave_reset_n;
  output           jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_3_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_3_avalon_jtag_slave_writedata;
  input            clk;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input            jtag_uart_3_avalon_jtag_slave_dataavailable;
  input            jtag_uart_3_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_3_avalon_jtag_slave_readdata;
  input            jtag_uart_3_avalon_jtag_slave_readyfordata;
  input            jtag_uart_3_avalon_jtag_slave_waitrequest;
  input            reset_n;

  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave;
  wire             cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave;
  wire             cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave;
  wire             cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave;
  wire             cpu_3_data_master_saved_grant_jtag_uart_3_avalon_jtag_slave;
  reg              d1_jtag_uart_3_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_3_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_3_avalon_jtag_slave_address;
  wire             jtag_uart_3_avalon_jtag_slave_allgrants;
  wire             jtag_uart_3_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_3_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_3_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_3_avalon_jtag_slave_arb_counter_enable;
  reg     [  2: 0] jtag_uart_3_avalon_jtag_slave_arb_share_counter;
  wire    [  2: 0] jtag_uart_3_avalon_jtag_slave_arb_share_counter_next_value;
  wire    [  2: 0] jtag_uart_3_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_3_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_3_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_3_avalon_jtag_slave_chipselect;
  wire             jtag_uart_3_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_3_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_3_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_3_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_3_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_3_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_3_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_3_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_3_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_3_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_3_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_3_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_3_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_3_avalon_jtag_slave_reset_n;
  reg              jtag_uart_3_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_3_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_3_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_3_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_3_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_3_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_3_avalon_jtag_slave_writedata;
  wire    [ 24: 0] shifted_address_to_jtag_uart_3_avalon_jtag_slave_from_cpu_3_data_master;
  wire             wait_for_jtag_uart_3_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_3_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_3_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave));
  //assign jtag_uart_3_avalon_jtag_slave_readdata_from_sa = jtag_uart_3_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_readdata_from_sa = jtag_uart_3_avalon_jtag_slave_readdata;

  assign cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave = ({cpu_3_data_master_address_to_slave[24 : 3] , 3'b0} == 25'h90) & (cpu_3_data_master_read | cpu_3_data_master_write);
  //assign jtag_uart_3_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_3_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_3_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_3_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_3_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_3_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_3_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_3_avalon_jtag_slave_waitrequest;

  //jtag_uart_3_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_3_avalon_jtag_slave_arb_share_set_values = 1;

  //jtag_uart_3_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_3_avalon_jtag_slave_non_bursting_master_requests = cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave;

  //jtag_uart_3_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_3_avalon_jtag_slave_any_bursting_master_saved_grant = 0;

  //jtag_uart_3_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_3_avalon_jtag_slave_firsttransfer ? (jtag_uart_3_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_3_avalon_jtag_slave_arb_share_counter ? (jtag_uart_3_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_3_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_3_avalon_jtag_slave_allgrants = |jtag_uart_3_avalon_jtag_slave_grant_vector;

  //jtag_uart_3_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_end_xfer = ~(jtag_uart_3_avalon_jtag_slave_waits_for_read | jtag_uart_3_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_3_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_3_avalon_jtag_slave = jtag_uart_3_avalon_jtag_slave_end_xfer & (~jtag_uart_3_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_3_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_3_avalon_jtag_slave & jtag_uart_3_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_3_avalon_jtag_slave & ~jtag_uart_3_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_3_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_3_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_3_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_3_avalon_jtag_slave_arb_share_counter <= jtag_uart_3_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_3_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_3_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_3_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_3_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_3_avalon_jtag_slave & ~jtag_uart_3_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_3_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_3_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //cpu_3/data_master jtag_uart_3/avalon_jtag_slave arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = jtag_uart_3_avalon_jtag_slave_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //jtag_uart_3_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_3_avalon_jtag_slave_arb_share_counter_next_value;

  //cpu_3/data_master jtag_uart_3/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = jtag_uart_3_avalon_jtag_slave_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //jtag_uart_3_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_any_continuerequest = 1;

  //cpu_3_data_master_continuerequest continued request, which is an e_assign
  assign cpu_3_data_master_continuerequest = 1;

  assign cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave = cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave & ~((cpu_3_data_master_read & ((cpu_3_data_master_latency_counter != 0) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))));
  //local readdatavalid cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave, which is an e_mux
  assign cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave = cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave & cpu_3_data_master_read & ~jtag_uart_3_avalon_jtag_slave_waits_for_read;

  //jtag_uart_3_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_3_avalon_jtag_slave_writedata = cpu_3_data_master_writedata;

  //master is always granted when requested
  assign cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave = cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave;

  //cpu_3/data_master saved-grant jtag_uart_3/avalon_jtag_slave, which is an e_assign
  assign cpu_3_data_master_saved_grant_jtag_uart_3_avalon_jtag_slave = cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart_3/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_3_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_3_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_3_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_3_avalon_jtag_slave_chipselect = cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave;
  //jtag_uart_3_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_firsttransfer = jtag_uart_3_avalon_jtag_slave_begins_xfer ? jtag_uart_3_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_3_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_3_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_3_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_3_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_3_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_3_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_3_avalon_jtag_slave_begins_xfer)
          jtag_uart_3_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_3_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_3_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_3_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_3_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_3_avalon_jtag_slave_read_n = ~(cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave & cpu_3_data_master_read);

  //~jtag_uart_3_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_3_avalon_jtag_slave_write_n = ~(cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave & cpu_3_data_master_write);

  assign shifted_address_to_jtag_uart_3_avalon_jtag_slave_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  //jtag_uart_3_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_3_avalon_jtag_slave_address = shifted_address_to_jtag_uart_3_avalon_jtag_slave_from_cpu_3_data_master >> 2;

  //d1_jtag_uart_3_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_3_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_3_avalon_jtag_slave_end_xfer <= jtag_uart_3_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_3_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_3_avalon_jtag_slave_waits_for_read = jtag_uart_3_avalon_jtag_slave_in_a_read_cycle & jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_3_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_in_a_read_cycle = cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave & cpu_3_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_3_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_3_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_3_avalon_jtag_slave_waits_for_write = jtag_uart_3_avalon_jtag_slave_in_a_write_cycle & jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_3_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_in_a_write_cycle = cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave & cpu_3_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_3_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_3_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_3_avalon_jtag_slave_irq_from_sa = jtag_uart_3_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_3_avalon_jtag_slave_irq_from_sa = jtag_uart_3_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart_3/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module keys_s1_arbitrator (
                            // inputs:
                             clk,
                             cpu_0_data_master_address_to_slave,
                             cpu_0_data_master_latency_counter,
                             cpu_0_data_master_read,
                             cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                             cpu_0_data_master_write,
                             cpu_0_data_master_writedata,
                             cpu_1_data_master_address_to_slave,
                             cpu_1_data_master_latency_counter,
                             cpu_1_data_master_read,
                             cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                             cpu_1_data_master_write,
                             cpu_1_data_master_writedata,
                             cpu_2_data_master_address_to_slave,
                             cpu_2_data_master_latency_counter,
                             cpu_2_data_master_read,
                             cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                             cpu_2_data_master_write,
                             cpu_2_data_master_writedata,
                             cpu_3_data_master_address_to_slave,
                             cpu_3_data_master_latency_counter,
                             cpu_3_data_master_read,
                             cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                             cpu_3_data_master_write,
                             cpu_3_data_master_writedata,
                             keys_s1_readdata,
                             reset_n,

                            // outputs:
                             cpu_0_data_master_granted_keys_s1,
                             cpu_0_data_master_qualified_request_keys_s1,
                             cpu_0_data_master_read_data_valid_keys_s1,
                             cpu_0_data_master_requests_keys_s1,
                             cpu_1_data_master_granted_keys_s1,
                             cpu_1_data_master_qualified_request_keys_s1,
                             cpu_1_data_master_read_data_valid_keys_s1,
                             cpu_1_data_master_requests_keys_s1,
                             cpu_2_data_master_granted_keys_s1,
                             cpu_2_data_master_qualified_request_keys_s1,
                             cpu_2_data_master_read_data_valid_keys_s1,
                             cpu_2_data_master_requests_keys_s1,
                             cpu_3_data_master_granted_keys_s1,
                             cpu_3_data_master_qualified_request_keys_s1,
                             cpu_3_data_master_read_data_valid_keys_s1,
                             cpu_3_data_master_requests_keys_s1,
                             d1_keys_s1_end_xfer,
                             keys_s1_address,
                             keys_s1_chipselect,
                             keys_s1_readdata_from_sa,
                             keys_s1_reset_n,
                             keys_s1_write_n,
                             keys_s1_writedata
                          )
;

  output           cpu_0_data_master_granted_keys_s1;
  output           cpu_0_data_master_qualified_request_keys_s1;
  output           cpu_0_data_master_read_data_valid_keys_s1;
  output           cpu_0_data_master_requests_keys_s1;
  output           cpu_1_data_master_granted_keys_s1;
  output           cpu_1_data_master_qualified_request_keys_s1;
  output           cpu_1_data_master_read_data_valid_keys_s1;
  output           cpu_1_data_master_requests_keys_s1;
  output           cpu_2_data_master_granted_keys_s1;
  output           cpu_2_data_master_qualified_request_keys_s1;
  output           cpu_2_data_master_read_data_valid_keys_s1;
  output           cpu_2_data_master_requests_keys_s1;
  output           cpu_3_data_master_granted_keys_s1;
  output           cpu_3_data_master_qualified_request_keys_s1;
  output           cpu_3_data_master_read_data_valid_keys_s1;
  output           cpu_3_data_master_requests_keys_s1;
  output           d1_keys_s1_end_xfer;
  output  [  1: 0] keys_s1_address;
  output           keys_s1_chipselect;
  output  [ 31: 0] keys_s1_readdata_from_sa;
  output           keys_s1_reset_n;
  output           keys_s1_write_n;
  output  [ 31: 0] keys_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 31: 0] keys_s1_readdata;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_keys_s1;
  wire             cpu_0_data_master_qualified_request_keys_s1;
  wire             cpu_0_data_master_read_data_valid_keys_s1;
  wire             cpu_0_data_master_requests_keys_s1;
  wire             cpu_0_data_master_saved_grant_keys_s1;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_keys_s1;
  wire             cpu_1_data_master_qualified_request_keys_s1;
  wire             cpu_1_data_master_read_data_valid_keys_s1;
  wire             cpu_1_data_master_requests_keys_s1;
  wire             cpu_1_data_master_saved_grant_keys_s1;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_keys_s1;
  wire             cpu_2_data_master_qualified_request_keys_s1;
  wire             cpu_2_data_master_read_data_valid_keys_s1;
  wire             cpu_2_data_master_requests_keys_s1;
  wire             cpu_2_data_master_saved_grant_keys_s1;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_keys_s1;
  wire             cpu_3_data_master_qualified_request_keys_s1;
  wire             cpu_3_data_master_read_data_valid_keys_s1;
  wire             cpu_3_data_master_requests_keys_s1;
  wire             cpu_3_data_master_saved_grant_keys_s1;
  reg              d1_keys_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_keys_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] keys_s1_address;
  wire             keys_s1_allgrants;
  wire             keys_s1_allow_new_arb_cycle;
  wire             keys_s1_any_bursting_master_saved_grant;
  wire             keys_s1_any_continuerequest;
  reg     [  3: 0] keys_s1_arb_addend;
  wire             keys_s1_arb_counter_enable;
  reg     [  2: 0] keys_s1_arb_share_counter;
  wire    [  2: 0] keys_s1_arb_share_counter_next_value;
  wire    [  2: 0] keys_s1_arb_share_set_values;
  wire    [  3: 0] keys_s1_arb_winner;
  wire             keys_s1_arbitration_holdoff_internal;
  wire             keys_s1_beginbursttransfer_internal;
  wire             keys_s1_begins_xfer;
  wire             keys_s1_chipselect;
  wire    [  7: 0] keys_s1_chosen_master_double_vector;
  wire    [  3: 0] keys_s1_chosen_master_rot_left;
  wire             keys_s1_end_xfer;
  wire             keys_s1_firsttransfer;
  wire    [  3: 0] keys_s1_grant_vector;
  wire             keys_s1_in_a_read_cycle;
  wire             keys_s1_in_a_write_cycle;
  wire    [  3: 0] keys_s1_master_qreq_vector;
  wire             keys_s1_non_bursting_master_requests;
  wire    [ 31: 0] keys_s1_readdata_from_sa;
  reg              keys_s1_reg_firsttransfer;
  wire             keys_s1_reset_n;
  reg     [  3: 0] keys_s1_saved_chosen_master_vector;
  reg              keys_s1_slavearbiterlockenable;
  wire             keys_s1_slavearbiterlockenable2;
  wire             keys_s1_unreg_firsttransfer;
  wire             keys_s1_waits_for_read;
  wire             keys_s1_waits_for_write;
  wire             keys_s1_write_n;
  wire    [ 31: 0] keys_s1_writedata;
  reg              last_cycle_cpu_0_data_master_granted_slave_keys_s1;
  reg              last_cycle_cpu_1_data_master_granted_slave_keys_s1;
  reg              last_cycle_cpu_2_data_master_granted_slave_keys_s1;
  reg              last_cycle_cpu_3_data_master_granted_slave_keys_s1;
  wire    [ 24: 0] shifted_address_to_keys_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_keys_s1_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_keys_s1_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_keys_s1_from_cpu_3_data_master;
  wire             wait_for_keys_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~keys_s1_end_xfer;
    end


  assign keys_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_keys_s1 | cpu_1_data_master_qualified_request_keys_s1 | cpu_2_data_master_qualified_request_keys_s1 | cpu_3_data_master_qualified_request_keys_s1));
  //assign keys_s1_readdata_from_sa = keys_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign keys_s1_readdata_from_sa = keys_s1_readdata;

  assign cpu_0_data_master_requests_keys_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h1903010) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //keys_s1_arb_share_counter set values, which is an e_mux
  assign keys_s1_arb_share_set_values = 1;

  //keys_s1_non_bursting_master_requests mux, which is an e_mux
  assign keys_s1_non_bursting_master_requests = cpu_0_data_master_requests_keys_s1 |
    cpu_1_data_master_requests_keys_s1 |
    cpu_2_data_master_requests_keys_s1 |
    cpu_3_data_master_requests_keys_s1 |
    cpu_0_data_master_requests_keys_s1 |
    cpu_1_data_master_requests_keys_s1 |
    cpu_2_data_master_requests_keys_s1 |
    cpu_3_data_master_requests_keys_s1 |
    cpu_0_data_master_requests_keys_s1 |
    cpu_1_data_master_requests_keys_s1 |
    cpu_2_data_master_requests_keys_s1 |
    cpu_3_data_master_requests_keys_s1 |
    cpu_0_data_master_requests_keys_s1 |
    cpu_1_data_master_requests_keys_s1 |
    cpu_2_data_master_requests_keys_s1 |
    cpu_3_data_master_requests_keys_s1;

  //keys_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign keys_s1_any_bursting_master_saved_grant = 0;

  //keys_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign keys_s1_arb_share_counter_next_value = keys_s1_firsttransfer ? (keys_s1_arb_share_set_values - 1) : |keys_s1_arb_share_counter ? (keys_s1_arb_share_counter - 1) : 0;

  //keys_s1_allgrants all slave grants, which is an e_mux
  assign keys_s1_allgrants = (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector) |
    (|keys_s1_grant_vector);

  //keys_s1_end_xfer assignment, which is an e_assign
  assign keys_s1_end_xfer = ~(keys_s1_waits_for_read | keys_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_keys_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_keys_s1 = keys_s1_end_xfer & (~keys_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //keys_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign keys_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_keys_s1 & keys_s1_allgrants) | (end_xfer_arb_share_counter_term_keys_s1 & ~keys_s1_non_bursting_master_requests);

  //keys_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          keys_s1_arb_share_counter <= 0;
      else if (keys_s1_arb_counter_enable)
          keys_s1_arb_share_counter <= keys_s1_arb_share_counter_next_value;
    end


  //keys_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          keys_s1_slavearbiterlockenable <= 0;
      else if ((|keys_s1_master_qreq_vector & end_xfer_arb_share_counter_term_keys_s1) | (end_xfer_arb_share_counter_term_keys_s1 & ~keys_s1_non_bursting_master_requests))
          keys_s1_slavearbiterlockenable <= |keys_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master keys/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = keys_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //keys_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign keys_s1_slavearbiterlockenable2 = |keys_s1_arb_share_counter_next_value;

  //cpu_0/data_master keys/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = keys_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_1/data_master keys/s1 arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = keys_s1_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master keys/s1 arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = keys_s1_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted keys/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_keys_s1 <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_keys_s1 <= cpu_1_data_master_saved_grant_keys_s1 ? 1 : (keys_s1_arbitration_holdoff_internal | ~cpu_1_data_master_requests_keys_s1) ? 0 : last_cycle_cpu_1_data_master_granted_slave_keys_s1;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_keys_s1 & cpu_1_data_master_requests_keys_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_keys_s1 & cpu_1_data_master_requests_keys_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_keys_s1 & cpu_1_data_master_requests_keys_s1);

  //keys_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign keys_s1_any_continuerequest = cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest;

  //cpu_2/data_master keys/s1 arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = keys_s1_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master keys/s1 arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = keys_s1_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted keys/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_keys_s1 <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_keys_s1 <= cpu_2_data_master_saved_grant_keys_s1 ? 1 : (keys_s1_arbitration_holdoff_internal | ~cpu_2_data_master_requests_keys_s1) ? 0 : last_cycle_cpu_2_data_master_granted_slave_keys_s1;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_keys_s1 & cpu_2_data_master_requests_keys_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_keys_s1 & cpu_2_data_master_requests_keys_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_keys_s1 & cpu_2_data_master_requests_keys_s1);

  //cpu_3/data_master keys/s1 arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = keys_s1_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master keys/s1 arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = keys_s1_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted keys/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_keys_s1 <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_keys_s1 <= cpu_3_data_master_saved_grant_keys_s1 ? 1 : (keys_s1_arbitration_holdoff_internal | ~cpu_3_data_master_requests_keys_s1) ? 0 : last_cycle_cpu_3_data_master_granted_slave_keys_s1;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_keys_s1 & cpu_3_data_master_requests_keys_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_keys_s1 & cpu_3_data_master_requests_keys_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_keys_s1 & cpu_3_data_master_requests_keys_s1);

  assign cpu_0_data_master_qualified_request_keys_s1 = cpu_0_data_master_requests_keys_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_keys_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_keys_s1 = cpu_0_data_master_granted_keys_s1 & cpu_0_data_master_read & ~keys_s1_waits_for_read;

  //keys_s1_writedata mux, which is an e_mux
  assign keys_s1_writedata = (cpu_0_data_master_granted_keys_s1)? cpu_0_data_master_writedata :
    (cpu_1_data_master_granted_keys_s1)? cpu_1_data_master_writedata :
    (cpu_2_data_master_granted_keys_s1)? cpu_2_data_master_writedata :
    cpu_3_data_master_writedata;

  assign cpu_1_data_master_requests_keys_s1 = ({cpu_1_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h1903010) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //cpu_0/data_master granted keys/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_keys_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_keys_s1 <= cpu_0_data_master_saved_grant_keys_s1 ? 1 : (keys_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_keys_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_keys_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_keys_s1 & cpu_0_data_master_requests_keys_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_keys_s1 & cpu_0_data_master_requests_keys_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_keys_s1 & cpu_0_data_master_requests_keys_s1);

  assign cpu_1_data_master_qualified_request_keys_s1 = cpu_1_data_master_requests_keys_s1 & ~((cpu_1_data_master_read & ((cpu_1_data_master_latency_counter != 0) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_1_data_master_read_data_valid_keys_s1, which is an e_mux
  assign cpu_1_data_master_read_data_valid_keys_s1 = cpu_1_data_master_granted_keys_s1 & cpu_1_data_master_read & ~keys_s1_waits_for_read;

  assign cpu_2_data_master_requests_keys_s1 = ({cpu_2_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h1903010) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_keys_s1 = cpu_2_data_master_requests_keys_s1 & ~((cpu_2_data_master_read & ((cpu_2_data_master_latency_counter != 0) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_2_data_master_read_data_valid_keys_s1, which is an e_mux
  assign cpu_2_data_master_read_data_valid_keys_s1 = cpu_2_data_master_granted_keys_s1 & cpu_2_data_master_read & ~keys_s1_waits_for_read;

  assign cpu_3_data_master_requests_keys_s1 = ({cpu_3_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h1903010) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_keys_s1 = cpu_3_data_master_requests_keys_s1 & ~((cpu_3_data_master_read & ((cpu_3_data_master_latency_counter != 0) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock);
  //local readdatavalid cpu_3_data_master_read_data_valid_keys_s1, which is an e_mux
  assign cpu_3_data_master_read_data_valid_keys_s1 = cpu_3_data_master_granted_keys_s1 & cpu_3_data_master_read & ~keys_s1_waits_for_read;

  //allow new arb cycle for keys/s1, which is an e_assign
  assign keys_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_3_data_master_arbiterlock;

  //cpu_3/data_master assignment into master qualified-requests vector for keys/s1, which is an e_assign
  assign keys_s1_master_qreq_vector[0] = cpu_3_data_master_qualified_request_keys_s1;

  //cpu_3/data_master grant keys/s1, which is an e_assign
  assign cpu_3_data_master_granted_keys_s1 = keys_s1_grant_vector[0];

  //cpu_3/data_master saved-grant keys/s1, which is an e_assign
  assign cpu_3_data_master_saved_grant_keys_s1 = keys_s1_arb_winner[0] && cpu_3_data_master_requests_keys_s1;

  //cpu_2/data_master assignment into master qualified-requests vector for keys/s1, which is an e_assign
  assign keys_s1_master_qreq_vector[1] = cpu_2_data_master_qualified_request_keys_s1;

  //cpu_2/data_master grant keys/s1, which is an e_assign
  assign cpu_2_data_master_granted_keys_s1 = keys_s1_grant_vector[1];

  //cpu_2/data_master saved-grant keys/s1, which is an e_assign
  assign cpu_2_data_master_saved_grant_keys_s1 = keys_s1_arb_winner[1] && cpu_2_data_master_requests_keys_s1;

  //cpu_1/data_master assignment into master qualified-requests vector for keys/s1, which is an e_assign
  assign keys_s1_master_qreq_vector[2] = cpu_1_data_master_qualified_request_keys_s1;

  //cpu_1/data_master grant keys/s1, which is an e_assign
  assign cpu_1_data_master_granted_keys_s1 = keys_s1_grant_vector[2];

  //cpu_1/data_master saved-grant keys/s1, which is an e_assign
  assign cpu_1_data_master_saved_grant_keys_s1 = keys_s1_arb_winner[2] && cpu_1_data_master_requests_keys_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for keys/s1, which is an e_assign
  assign keys_s1_master_qreq_vector[3] = cpu_0_data_master_qualified_request_keys_s1;

  //cpu_0/data_master grant keys/s1, which is an e_assign
  assign cpu_0_data_master_granted_keys_s1 = keys_s1_grant_vector[3];

  //cpu_0/data_master saved-grant keys/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_keys_s1 = keys_s1_arb_winner[3] && cpu_0_data_master_requests_keys_s1;

  //keys/s1 chosen-master double-vector, which is an e_assign
  assign keys_s1_chosen_master_double_vector = {keys_s1_master_qreq_vector, keys_s1_master_qreq_vector} & ({~keys_s1_master_qreq_vector, ~keys_s1_master_qreq_vector} + keys_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign keys_s1_arb_winner = (keys_s1_allow_new_arb_cycle & | keys_s1_grant_vector) ? keys_s1_grant_vector : keys_s1_saved_chosen_master_vector;

  //saved keys_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          keys_s1_saved_chosen_master_vector <= 0;
      else if (keys_s1_allow_new_arb_cycle)
          keys_s1_saved_chosen_master_vector <= |keys_s1_grant_vector ? keys_s1_grant_vector : keys_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign keys_s1_grant_vector = {(keys_s1_chosen_master_double_vector[3] | keys_s1_chosen_master_double_vector[7]),
    (keys_s1_chosen_master_double_vector[2] | keys_s1_chosen_master_double_vector[6]),
    (keys_s1_chosen_master_double_vector[1] | keys_s1_chosen_master_double_vector[5]),
    (keys_s1_chosen_master_double_vector[0] | keys_s1_chosen_master_double_vector[4])};

  //keys/s1 chosen master rotated left, which is an e_assign
  assign keys_s1_chosen_master_rot_left = (keys_s1_arb_winner << 1) ? (keys_s1_arb_winner << 1) : 1;

  //keys/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          keys_s1_arb_addend <= 1;
      else if (|keys_s1_grant_vector)
          keys_s1_arb_addend <= keys_s1_end_xfer? keys_s1_chosen_master_rot_left : keys_s1_grant_vector;
    end


  //keys_s1_reset_n assignment, which is an e_assign
  assign keys_s1_reset_n = reset_n;

  assign keys_s1_chipselect = cpu_0_data_master_granted_keys_s1 | cpu_1_data_master_granted_keys_s1 | cpu_2_data_master_granted_keys_s1 | cpu_3_data_master_granted_keys_s1;
  //keys_s1_firsttransfer first transaction, which is an e_assign
  assign keys_s1_firsttransfer = keys_s1_begins_xfer ? keys_s1_unreg_firsttransfer : keys_s1_reg_firsttransfer;

  //keys_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign keys_s1_unreg_firsttransfer = ~(keys_s1_slavearbiterlockenable & keys_s1_any_continuerequest);

  //keys_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          keys_s1_reg_firsttransfer <= 1'b1;
      else if (keys_s1_begins_xfer)
          keys_s1_reg_firsttransfer <= keys_s1_unreg_firsttransfer;
    end


  //keys_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign keys_s1_beginbursttransfer_internal = keys_s1_begins_xfer;

  //keys_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign keys_s1_arbitration_holdoff_internal = keys_s1_begins_xfer & keys_s1_firsttransfer;

  //~keys_s1_write_n assignment, which is an e_mux
  assign keys_s1_write_n = ~((cpu_0_data_master_granted_keys_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_keys_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_keys_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_keys_s1 & cpu_3_data_master_write));

  assign shifted_address_to_keys_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //keys_s1_address mux, which is an e_mux
  assign keys_s1_address = (cpu_0_data_master_granted_keys_s1)? (shifted_address_to_keys_s1_from_cpu_0_data_master >> 2) :
    (cpu_1_data_master_granted_keys_s1)? (shifted_address_to_keys_s1_from_cpu_1_data_master >> 2) :
    (cpu_2_data_master_granted_keys_s1)? (shifted_address_to_keys_s1_from_cpu_2_data_master >> 2) :
    (shifted_address_to_keys_s1_from_cpu_3_data_master >> 2);

  assign shifted_address_to_keys_s1_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_keys_s1_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_keys_s1_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  //d1_keys_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_keys_s1_end_xfer <= 1;
      else 
        d1_keys_s1_end_xfer <= keys_s1_end_xfer;
    end


  //keys_s1_waits_for_read in a cycle, which is an e_mux
  assign keys_s1_waits_for_read = keys_s1_in_a_read_cycle & keys_s1_begins_xfer;

  //keys_s1_in_a_read_cycle assignment, which is an e_assign
  assign keys_s1_in_a_read_cycle = (cpu_0_data_master_granted_keys_s1 & cpu_0_data_master_read) | (cpu_1_data_master_granted_keys_s1 & cpu_1_data_master_read) | (cpu_2_data_master_granted_keys_s1 & cpu_2_data_master_read) | (cpu_3_data_master_granted_keys_s1 & cpu_3_data_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = keys_s1_in_a_read_cycle;

  //keys_s1_waits_for_write in a cycle, which is an e_mux
  assign keys_s1_waits_for_write = keys_s1_in_a_write_cycle & 0;

  //keys_s1_in_a_write_cycle assignment, which is an e_assign
  assign keys_s1_in_a_write_cycle = (cpu_0_data_master_granted_keys_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_keys_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_keys_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_keys_s1 & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = keys_s1_in_a_write_cycle;

  assign wait_for_keys_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //keys/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_keys_s1 + cpu_1_data_master_granted_keys_s1 + cpu_2_data_master_granted_keys_s1 + cpu_3_data_master_granted_keys_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_keys_s1 + cpu_1_data_master_saved_grant_keys_s1 + cpu_2_data_master_saved_grant_keys_s1 + cpu_3_data_master_saved_grant_keys_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module mailbox_0_s1_arbitrator (
                                 // inputs:
                                  clk,
                                  cpu_0_data_master_address_to_slave,
                                  cpu_0_data_master_latency_counter,
                                  cpu_0_data_master_read,
                                  cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_0_data_master_write,
                                  cpu_0_data_master_writedata,
                                  cpu_1_data_master_address_to_slave,
                                  cpu_1_data_master_latency_counter,
                                  cpu_1_data_master_read,
                                  cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_1_data_master_write,
                                  cpu_1_data_master_writedata,
                                  cpu_2_data_master_address_to_slave,
                                  cpu_2_data_master_latency_counter,
                                  cpu_2_data_master_read,
                                  cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_2_data_master_write,
                                  cpu_2_data_master_writedata,
                                  cpu_3_data_master_address_to_slave,
                                  cpu_3_data_master_latency_counter,
                                  cpu_3_data_master_read,
                                  cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_3_data_master_write,
                                  cpu_3_data_master_writedata,
                                  mailbox_0_s1_readdata,
                                  reset_n,

                                 // outputs:
                                  cpu_0_data_master_granted_mailbox_0_s1,
                                  cpu_0_data_master_qualified_request_mailbox_0_s1,
                                  cpu_0_data_master_read_data_valid_mailbox_0_s1,
                                  cpu_0_data_master_requests_mailbox_0_s1,
                                  cpu_1_data_master_granted_mailbox_0_s1,
                                  cpu_1_data_master_qualified_request_mailbox_0_s1,
                                  cpu_1_data_master_read_data_valid_mailbox_0_s1,
                                  cpu_1_data_master_requests_mailbox_0_s1,
                                  cpu_2_data_master_granted_mailbox_0_s1,
                                  cpu_2_data_master_qualified_request_mailbox_0_s1,
                                  cpu_2_data_master_read_data_valid_mailbox_0_s1,
                                  cpu_2_data_master_requests_mailbox_0_s1,
                                  cpu_3_data_master_granted_mailbox_0_s1,
                                  cpu_3_data_master_qualified_request_mailbox_0_s1,
                                  cpu_3_data_master_read_data_valid_mailbox_0_s1,
                                  cpu_3_data_master_requests_mailbox_0_s1,
                                  d1_mailbox_0_s1_end_xfer,
                                  mailbox_0_s1_address,
                                  mailbox_0_s1_chipselect,
                                  mailbox_0_s1_read,
                                  mailbox_0_s1_readdata_from_sa,
                                  mailbox_0_s1_reset_n,
                                  mailbox_0_s1_write,
                                  mailbox_0_s1_writedata
                               )
;

  output           cpu_0_data_master_granted_mailbox_0_s1;
  output           cpu_0_data_master_qualified_request_mailbox_0_s1;
  output           cpu_0_data_master_read_data_valid_mailbox_0_s1;
  output           cpu_0_data_master_requests_mailbox_0_s1;
  output           cpu_1_data_master_granted_mailbox_0_s1;
  output           cpu_1_data_master_qualified_request_mailbox_0_s1;
  output           cpu_1_data_master_read_data_valid_mailbox_0_s1;
  output           cpu_1_data_master_requests_mailbox_0_s1;
  output           cpu_2_data_master_granted_mailbox_0_s1;
  output           cpu_2_data_master_qualified_request_mailbox_0_s1;
  output           cpu_2_data_master_read_data_valid_mailbox_0_s1;
  output           cpu_2_data_master_requests_mailbox_0_s1;
  output           cpu_3_data_master_granted_mailbox_0_s1;
  output           cpu_3_data_master_qualified_request_mailbox_0_s1;
  output           cpu_3_data_master_read_data_valid_mailbox_0_s1;
  output           cpu_3_data_master_requests_mailbox_0_s1;
  output           d1_mailbox_0_s1_end_xfer;
  output  [  1: 0] mailbox_0_s1_address;
  output           mailbox_0_s1_chipselect;
  output           mailbox_0_s1_read;
  output  [ 31: 0] mailbox_0_s1_readdata_from_sa;
  output           mailbox_0_s1_reset_n;
  output           mailbox_0_s1_write;
  output  [ 31: 0] mailbox_0_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 31: 0] mailbox_0_s1_readdata;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_mailbox_0_s1;
  wire             cpu_0_data_master_qualified_request_mailbox_0_s1;
  wire             cpu_0_data_master_read_data_valid_mailbox_0_s1;
  wire             cpu_0_data_master_requests_mailbox_0_s1;
  wire             cpu_0_data_master_saved_grant_mailbox_0_s1;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_mailbox_0_s1;
  wire             cpu_1_data_master_qualified_request_mailbox_0_s1;
  wire             cpu_1_data_master_read_data_valid_mailbox_0_s1;
  wire             cpu_1_data_master_requests_mailbox_0_s1;
  wire             cpu_1_data_master_saved_grant_mailbox_0_s1;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_mailbox_0_s1;
  wire             cpu_2_data_master_qualified_request_mailbox_0_s1;
  wire             cpu_2_data_master_read_data_valid_mailbox_0_s1;
  wire             cpu_2_data_master_requests_mailbox_0_s1;
  wire             cpu_2_data_master_saved_grant_mailbox_0_s1;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_mailbox_0_s1;
  wire             cpu_3_data_master_qualified_request_mailbox_0_s1;
  wire             cpu_3_data_master_read_data_valid_mailbox_0_s1;
  wire             cpu_3_data_master_requests_mailbox_0_s1;
  wire             cpu_3_data_master_saved_grant_mailbox_0_s1;
  reg              d1_mailbox_0_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_mailbox_0_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_mailbox_0_s1;
  reg              last_cycle_cpu_1_data_master_granted_slave_mailbox_0_s1;
  reg              last_cycle_cpu_2_data_master_granted_slave_mailbox_0_s1;
  reg              last_cycle_cpu_3_data_master_granted_slave_mailbox_0_s1;
  wire    [  1: 0] mailbox_0_s1_address;
  wire             mailbox_0_s1_allgrants;
  wire             mailbox_0_s1_allow_new_arb_cycle;
  wire             mailbox_0_s1_any_bursting_master_saved_grant;
  wire             mailbox_0_s1_any_continuerequest;
  reg     [  3: 0] mailbox_0_s1_arb_addend;
  wire             mailbox_0_s1_arb_counter_enable;
  reg     [  2: 0] mailbox_0_s1_arb_share_counter;
  wire    [  2: 0] mailbox_0_s1_arb_share_counter_next_value;
  wire    [  2: 0] mailbox_0_s1_arb_share_set_values;
  wire    [  3: 0] mailbox_0_s1_arb_winner;
  wire             mailbox_0_s1_arbitration_holdoff_internal;
  wire             mailbox_0_s1_beginbursttransfer_internal;
  wire             mailbox_0_s1_begins_xfer;
  wire             mailbox_0_s1_chipselect;
  wire    [  7: 0] mailbox_0_s1_chosen_master_double_vector;
  wire    [  3: 0] mailbox_0_s1_chosen_master_rot_left;
  wire             mailbox_0_s1_end_xfer;
  wire             mailbox_0_s1_firsttransfer;
  wire    [  3: 0] mailbox_0_s1_grant_vector;
  wire             mailbox_0_s1_in_a_read_cycle;
  wire             mailbox_0_s1_in_a_write_cycle;
  wire    [  3: 0] mailbox_0_s1_master_qreq_vector;
  wire             mailbox_0_s1_non_bursting_master_requests;
  wire             mailbox_0_s1_read;
  wire    [ 31: 0] mailbox_0_s1_readdata_from_sa;
  reg              mailbox_0_s1_reg_firsttransfer;
  wire             mailbox_0_s1_reset_n;
  reg     [  3: 0] mailbox_0_s1_saved_chosen_master_vector;
  reg              mailbox_0_s1_slavearbiterlockenable;
  wire             mailbox_0_s1_slavearbiterlockenable2;
  wire             mailbox_0_s1_unreg_firsttransfer;
  wire             mailbox_0_s1_waits_for_read;
  wire             mailbox_0_s1_waits_for_write;
  wire             mailbox_0_s1_write;
  wire    [ 31: 0] mailbox_0_s1_writedata;
  wire    [ 24: 0] shifted_address_to_mailbox_0_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_0_s1_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_0_s1_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_0_s1_from_cpu_3_data_master;
  wire             wait_for_mailbox_0_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~mailbox_0_s1_end_xfer;
    end


  assign mailbox_0_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_mailbox_0_s1 | cpu_1_data_master_qualified_request_mailbox_0_s1 | cpu_2_data_master_qualified_request_mailbox_0_s1 | cpu_3_data_master_qualified_request_mailbox_0_s1));
  //assign mailbox_0_s1_readdata_from_sa = mailbox_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign mailbox_0_s1_readdata_from_sa = mailbox_0_s1_readdata;

  assign cpu_0_data_master_requests_mailbox_0_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h40) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //mailbox_0_s1_arb_share_counter set values, which is an e_mux
  assign mailbox_0_s1_arb_share_set_values = 1;

  //mailbox_0_s1_non_bursting_master_requests mux, which is an e_mux
  assign mailbox_0_s1_non_bursting_master_requests = cpu_0_data_master_requests_mailbox_0_s1 |
    cpu_1_data_master_requests_mailbox_0_s1 |
    cpu_2_data_master_requests_mailbox_0_s1 |
    cpu_3_data_master_requests_mailbox_0_s1 |
    cpu_0_data_master_requests_mailbox_0_s1 |
    cpu_1_data_master_requests_mailbox_0_s1 |
    cpu_2_data_master_requests_mailbox_0_s1 |
    cpu_3_data_master_requests_mailbox_0_s1 |
    cpu_0_data_master_requests_mailbox_0_s1 |
    cpu_1_data_master_requests_mailbox_0_s1 |
    cpu_2_data_master_requests_mailbox_0_s1 |
    cpu_3_data_master_requests_mailbox_0_s1 |
    cpu_0_data_master_requests_mailbox_0_s1 |
    cpu_1_data_master_requests_mailbox_0_s1 |
    cpu_2_data_master_requests_mailbox_0_s1 |
    cpu_3_data_master_requests_mailbox_0_s1;

  //mailbox_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign mailbox_0_s1_any_bursting_master_saved_grant = 0;

  //mailbox_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign mailbox_0_s1_arb_share_counter_next_value = mailbox_0_s1_firsttransfer ? (mailbox_0_s1_arb_share_set_values - 1) : |mailbox_0_s1_arb_share_counter ? (mailbox_0_s1_arb_share_counter - 1) : 0;

  //mailbox_0_s1_allgrants all slave grants, which is an e_mux
  assign mailbox_0_s1_allgrants = (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector) |
    (|mailbox_0_s1_grant_vector);

  //mailbox_0_s1_end_xfer assignment, which is an e_assign
  assign mailbox_0_s1_end_xfer = ~(mailbox_0_s1_waits_for_read | mailbox_0_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_mailbox_0_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_mailbox_0_s1 = mailbox_0_s1_end_xfer & (~mailbox_0_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //mailbox_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign mailbox_0_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_mailbox_0_s1 & mailbox_0_s1_allgrants) | (end_xfer_arb_share_counter_term_mailbox_0_s1 & ~mailbox_0_s1_non_bursting_master_requests);

  //mailbox_0_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_0_s1_arb_share_counter <= 0;
      else if (mailbox_0_s1_arb_counter_enable)
          mailbox_0_s1_arb_share_counter <= mailbox_0_s1_arb_share_counter_next_value;
    end


  //mailbox_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_0_s1_slavearbiterlockenable <= 0;
      else if ((|mailbox_0_s1_master_qreq_vector & end_xfer_arb_share_counter_term_mailbox_0_s1) | (end_xfer_arb_share_counter_term_mailbox_0_s1 & ~mailbox_0_s1_non_bursting_master_requests))
          mailbox_0_s1_slavearbiterlockenable <= |mailbox_0_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master mailbox_0/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = mailbox_0_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //mailbox_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign mailbox_0_s1_slavearbiterlockenable2 = |mailbox_0_s1_arb_share_counter_next_value;

  //cpu_0/data_master mailbox_0/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = mailbox_0_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_1/data_master mailbox_0/s1 arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = mailbox_0_s1_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master mailbox_0/s1 arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = mailbox_0_s1_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted mailbox_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_mailbox_0_s1 <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_mailbox_0_s1 <= cpu_1_data_master_saved_grant_mailbox_0_s1 ? 1 : (mailbox_0_s1_arbitration_holdoff_internal | ~cpu_1_data_master_requests_mailbox_0_s1) ? 0 : last_cycle_cpu_1_data_master_granted_slave_mailbox_0_s1;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_mailbox_0_s1 & cpu_1_data_master_requests_mailbox_0_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_mailbox_0_s1 & cpu_1_data_master_requests_mailbox_0_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_mailbox_0_s1 & cpu_1_data_master_requests_mailbox_0_s1);

  //mailbox_0_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign mailbox_0_s1_any_continuerequest = cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest;

  //cpu_2/data_master mailbox_0/s1 arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = mailbox_0_s1_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master mailbox_0/s1 arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = mailbox_0_s1_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted mailbox_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_mailbox_0_s1 <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_mailbox_0_s1 <= cpu_2_data_master_saved_grant_mailbox_0_s1 ? 1 : (mailbox_0_s1_arbitration_holdoff_internal | ~cpu_2_data_master_requests_mailbox_0_s1) ? 0 : last_cycle_cpu_2_data_master_granted_slave_mailbox_0_s1;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_mailbox_0_s1 & cpu_2_data_master_requests_mailbox_0_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_mailbox_0_s1 & cpu_2_data_master_requests_mailbox_0_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_mailbox_0_s1 & cpu_2_data_master_requests_mailbox_0_s1);

  //cpu_3/data_master mailbox_0/s1 arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = mailbox_0_s1_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master mailbox_0/s1 arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = mailbox_0_s1_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted mailbox_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_mailbox_0_s1 <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_mailbox_0_s1 <= cpu_3_data_master_saved_grant_mailbox_0_s1 ? 1 : (mailbox_0_s1_arbitration_holdoff_internal | ~cpu_3_data_master_requests_mailbox_0_s1) ? 0 : last_cycle_cpu_3_data_master_granted_slave_mailbox_0_s1;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_mailbox_0_s1 & cpu_3_data_master_requests_mailbox_0_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_mailbox_0_s1 & cpu_3_data_master_requests_mailbox_0_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_mailbox_0_s1 & cpu_3_data_master_requests_mailbox_0_s1);

  assign cpu_0_data_master_qualified_request_mailbox_0_s1 = cpu_0_data_master_requests_mailbox_0_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_mailbox_0_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_mailbox_0_s1 = cpu_0_data_master_granted_mailbox_0_s1 & cpu_0_data_master_read & ~mailbox_0_s1_waits_for_read;

  //mailbox_0_s1_writedata mux, which is an e_mux
  assign mailbox_0_s1_writedata = (cpu_0_data_master_granted_mailbox_0_s1)? cpu_0_data_master_writedata :
    (cpu_1_data_master_granted_mailbox_0_s1)? cpu_1_data_master_writedata :
    (cpu_2_data_master_granted_mailbox_0_s1)? cpu_2_data_master_writedata :
    cpu_3_data_master_writedata;

  assign cpu_1_data_master_requests_mailbox_0_s1 = ({cpu_1_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h40) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //cpu_0/data_master granted mailbox_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_mailbox_0_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_mailbox_0_s1 <= cpu_0_data_master_saved_grant_mailbox_0_s1 ? 1 : (mailbox_0_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_mailbox_0_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_mailbox_0_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_mailbox_0_s1 & cpu_0_data_master_requests_mailbox_0_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_mailbox_0_s1 & cpu_0_data_master_requests_mailbox_0_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_mailbox_0_s1 & cpu_0_data_master_requests_mailbox_0_s1);

  assign cpu_1_data_master_qualified_request_mailbox_0_s1 = cpu_1_data_master_requests_mailbox_0_s1 & ~((cpu_1_data_master_read & ((cpu_1_data_master_latency_counter != 0) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_1_data_master_read_data_valid_mailbox_0_s1, which is an e_mux
  assign cpu_1_data_master_read_data_valid_mailbox_0_s1 = cpu_1_data_master_granted_mailbox_0_s1 & cpu_1_data_master_read & ~mailbox_0_s1_waits_for_read;

  assign cpu_2_data_master_requests_mailbox_0_s1 = ({cpu_2_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h40) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_mailbox_0_s1 = cpu_2_data_master_requests_mailbox_0_s1 & ~((cpu_2_data_master_read & ((cpu_2_data_master_latency_counter != 0) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_2_data_master_read_data_valid_mailbox_0_s1, which is an e_mux
  assign cpu_2_data_master_read_data_valid_mailbox_0_s1 = cpu_2_data_master_granted_mailbox_0_s1 & cpu_2_data_master_read & ~mailbox_0_s1_waits_for_read;

  assign cpu_3_data_master_requests_mailbox_0_s1 = ({cpu_3_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h40) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_mailbox_0_s1 = cpu_3_data_master_requests_mailbox_0_s1 & ~((cpu_3_data_master_read & ((cpu_3_data_master_latency_counter != 0) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock);
  //local readdatavalid cpu_3_data_master_read_data_valid_mailbox_0_s1, which is an e_mux
  assign cpu_3_data_master_read_data_valid_mailbox_0_s1 = cpu_3_data_master_granted_mailbox_0_s1 & cpu_3_data_master_read & ~mailbox_0_s1_waits_for_read;

  //allow new arb cycle for mailbox_0/s1, which is an e_assign
  assign mailbox_0_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_3_data_master_arbiterlock;

  //cpu_3/data_master assignment into master qualified-requests vector for mailbox_0/s1, which is an e_assign
  assign mailbox_0_s1_master_qreq_vector[0] = cpu_3_data_master_qualified_request_mailbox_0_s1;

  //cpu_3/data_master grant mailbox_0/s1, which is an e_assign
  assign cpu_3_data_master_granted_mailbox_0_s1 = mailbox_0_s1_grant_vector[0];

  //cpu_3/data_master saved-grant mailbox_0/s1, which is an e_assign
  assign cpu_3_data_master_saved_grant_mailbox_0_s1 = mailbox_0_s1_arb_winner[0] && cpu_3_data_master_requests_mailbox_0_s1;

  //cpu_2/data_master assignment into master qualified-requests vector for mailbox_0/s1, which is an e_assign
  assign mailbox_0_s1_master_qreq_vector[1] = cpu_2_data_master_qualified_request_mailbox_0_s1;

  //cpu_2/data_master grant mailbox_0/s1, which is an e_assign
  assign cpu_2_data_master_granted_mailbox_0_s1 = mailbox_0_s1_grant_vector[1];

  //cpu_2/data_master saved-grant mailbox_0/s1, which is an e_assign
  assign cpu_2_data_master_saved_grant_mailbox_0_s1 = mailbox_0_s1_arb_winner[1] && cpu_2_data_master_requests_mailbox_0_s1;

  //cpu_1/data_master assignment into master qualified-requests vector for mailbox_0/s1, which is an e_assign
  assign mailbox_0_s1_master_qreq_vector[2] = cpu_1_data_master_qualified_request_mailbox_0_s1;

  //cpu_1/data_master grant mailbox_0/s1, which is an e_assign
  assign cpu_1_data_master_granted_mailbox_0_s1 = mailbox_0_s1_grant_vector[2];

  //cpu_1/data_master saved-grant mailbox_0/s1, which is an e_assign
  assign cpu_1_data_master_saved_grant_mailbox_0_s1 = mailbox_0_s1_arb_winner[2] && cpu_1_data_master_requests_mailbox_0_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for mailbox_0/s1, which is an e_assign
  assign mailbox_0_s1_master_qreq_vector[3] = cpu_0_data_master_qualified_request_mailbox_0_s1;

  //cpu_0/data_master grant mailbox_0/s1, which is an e_assign
  assign cpu_0_data_master_granted_mailbox_0_s1 = mailbox_0_s1_grant_vector[3];

  //cpu_0/data_master saved-grant mailbox_0/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_mailbox_0_s1 = mailbox_0_s1_arb_winner[3] && cpu_0_data_master_requests_mailbox_0_s1;

  //mailbox_0/s1 chosen-master double-vector, which is an e_assign
  assign mailbox_0_s1_chosen_master_double_vector = {mailbox_0_s1_master_qreq_vector, mailbox_0_s1_master_qreq_vector} & ({~mailbox_0_s1_master_qreq_vector, ~mailbox_0_s1_master_qreq_vector} + mailbox_0_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign mailbox_0_s1_arb_winner = (mailbox_0_s1_allow_new_arb_cycle & | mailbox_0_s1_grant_vector) ? mailbox_0_s1_grant_vector : mailbox_0_s1_saved_chosen_master_vector;

  //saved mailbox_0_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_0_s1_saved_chosen_master_vector <= 0;
      else if (mailbox_0_s1_allow_new_arb_cycle)
          mailbox_0_s1_saved_chosen_master_vector <= |mailbox_0_s1_grant_vector ? mailbox_0_s1_grant_vector : mailbox_0_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign mailbox_0_s1_grant_vector = {(mailbox_0_s1_chosen_master_double_vector[3] | mailbox_0_s1_chosen_master_double_vector[7]),
    (mailbox_0_s1_chosen_master_double_vector[2] | mailbox_0_s1_chosen_master_double_vector[6]),
    (mailbox_0_s1_chosen_master_double_vector[1] | mailbox_0_s1_chosen_master_double_vector[5]),
    (mailbox_0_s1_chosen_master_double_vector[0] | mailbox_0_s1_chosen_master_double_vector[4])};

  //mailbox_0/s1 chosen master rotated left, which is an e_assign
  assign mailbox_0_s1_chosen_master_rot_left = (mailbox_0_s1_arb_winner << 1) ? (mailbox_0_s1_arb_winner << 1) : 1;

  //mailbox_0/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_0_s1_arb_addend <= 1;
      else if (|mailbox_0_s1_grant_vector)
          mailbox_0_s1_arb_addend <= mailbox_0_s1_end_xfer? mailbox_0_s1_chosen_master_rot_left : mailbox_0_s1_grant_vector;
    end


  //mailbox_0_s1_reset_n assignment, which is an e_assign
  assign mailbox_0_s1_reset_n = reset_n;

  assign mailbox_0_s1_chipselect = cpu_0_data_master_granted_mailbox_0_s1 | cpu_1_data_master_granted_mailbox_0_s1 | cpu_2_data_master_granted_mailbox_0_s1 | cpu_3_data_master_granted_mailbox_0_s1;
  //mailbox_0_s1_firsttransfer first transaction, which is an e_assign
  assign mailbox_0_s1_firsttransfer = mailbox_0_s1_begins_xfer ? mailbox_0_s1_unreg_firsttransfer : mailbox_0_s1_reg_firsttransfer;

  //mailbox_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign mailbox_0_s1_unreg_firsttransfer = ~(mailbox_0_s1_slavearbiterlockenable & mailbox_0_s1_any_continuerequest);

  //mailbox_0_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_0_s1_reg_firsttransfer <= 1'b1;
      else if (mailbox_0_s1_begins_xfer)
          mailbox_0_s1_reg_firsttransfer <= mailbox_0_s1_unreg_firsttransfer;
    end


  //mailbox_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign mailbox_0_s1_beginbursttransfer_internal = mailbox_0_s1_begins_xfer;

  //mailbox_0_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign mailbox_0_s1_arbitration_holdoff_internal = mailbox_0_s1_begins_xfer & mailbox_0_s1_firsttransfer;

  //mailbox_0_s1_read assignment, which is an e_mux
  assign mailbox_0_s1_read = (cpu_0_data_master_granted_mailbox_0_s1 & cpu_0_data_master_read) | (cpu_1_data_master_granted_mailbox_0_s1 & cpu_1_data_master_read) | (cpu_2_data_master_granted_mailbox_0_s1 & cpu_2_data_master_read) | (cpu_3_data_master_granted_mailbox_0_s1 & cpu_3_data_master_read);

  //mailbox_0_s1_write assignment, which is an e_mux
  assign mailbox_0_s1_write = (cpu_0_data_master_granted_mailbox_0_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_mailbox_0_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_mailbox_0_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_mailbox_0_s1 & cpu_3_data_master_write);

  assign shifted_address_to_mailbox_0_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //mailbox_0_s1_address mux, which is an e_mux
  assign mailbox_0_s1_address = (cpu_0_data_master_granted_mailbox_0_s1)? (shifted_address_to_mailbox_0_s1_from_cpu_0_data_master >> 2) :
    (cpu_1_data_master_granted_mailbox_0_s1)? (shifted_address_to_mailbox_0_s1_from_cpu_1_data_master >> 2) :
    (cpu_2_data_master_granted_mailbox_0_s1)? (shifted_address_to_mailbox_0_s1_from_cpu_2_data_master >> 2) :
    (shifted_address_to_mailbox_0_s1_from_cpu_3_data_master >> 2);

  assign shifted_address_to_mailbox_0_s1_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_mailbox_0_s1_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_mailbox_0_s1_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  //d1_mailbox_0_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_mailbox_0_s1_end_xfer <= 1;
      else 
        d1_mailbox_0_s1_end_xfer <= mailbox_0_s1_end_xfer;
    end


  //mailbox_0_s1_waits_for_read in a cycle, which is an e_mux
  assign mailbox_0_s1_waits_for_read = mailbox_0_s1_in_a_read_cycle & mailbox_0_s1_begins_xfer;

  //mailbox_0_s1_in_a_read_cycle assignment, which is an e_assign
  assign mailbox_0_s1_in_a_read_cycle = (cpu_0_data_master_granted_mailbox_0_s1 & cpu_0_data_master_read) | (cpu_1_data_master_granted_mailbox_0_s1 & cpu_1_data_master_read) | (cpu_2_data_master_granted_mailbox_0_s1 & cpu_2_data_master_read) | (cpu_3_data_master_granted_mailbox_0_s1 & cpu_3_data_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = mailbox_0_s1_in_a_read_cycle;

  //mailbox_0_s1_waits_for_write in a cycle, which is an e_mux
  assign mailbox_0_s1_waits_for_write = mailbox_0_s1_in_a_write_cycle & 0;

  //mailbox_0_s1_in_a_write_cycle assignment, which is an e_assign
  assign mailbox_0_s1_in_a_write_cycle = (cpu_0_data_master_granted_mailbox_0_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_mailbox_0_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_mailbox_0_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_mailbox_0_s1 & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = mailbox_0_s1_in_a_write_cycle;

  assign wait_for_mailbox_0_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //mailbox_0/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_mailbox_0_s1 + cpu_1_data_master_granted_mailbox_0_s1 + cpu_2_data_master_granted_mailbox_0_s1 + cpu_3_data_master_granted_mailbox_0_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_mailbox_0_s1 + cpu_1_data_master_saved_grant_mailbox_0_s1 + cpu_2_data_master_saved_grant_mailbox_0_s1 + cpu_3_data_master_saved_grant_mailbox_0_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module mailbox_1_s1_arbitrator (
                                 // inputs:
                                  clk,
                                  cpu_0_data_master_address_to_slave,
                                  cpu_0_data_master_latency_counter,
                                  cpu_0_data_master_read,
                                  cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_0_data_master_write,
                                  cpu_0_data_master_writedata,
                                  cpu_1_data_master_address_to_slave,
                                  cpu_1_data_master_latency_counter,
                                  cpu_1_data_master_read,
                                  cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_1_data_master_write,
                                  cpu_1_data_master_writedata,
                                  cpu_2_data_master_address_to_slave,
                                  cpu_2_data_master_latency_counter,
                                  cpu_2_data_master_read,
                                  cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_2_data_master_write,
                                  cpu_2_data_master_writedata,
                                  cpu_3_data_master_address_to_slave,
                                  cpu_3_data_master_latency_counter,
                                  cpu_3_data_master_read,
                                  cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_3_data_master_write,
                                  cpu_3_data_master_writedata,
                                  mailbox_1_s1_readdata,
                                  reset_n,

                                 // outputs:
                                  cpu_0_data_master_granted_mailbox_1_s1,
                                  cpu_0_data_master_qualified_request_mailbox_1_s1,
                                  cpu_0_data_master_read_data_valid_mailbox_1_s1,
                                  cpu_0_data_master_requests_mailbox_1_s1,
                                  cpu_1_data_master_granted_mailbox_1_s1,
                                  cpu_1_data_master_qualified_request_mailbox_1_s1,
                                  cpu_1_data_master_read_data_valid_mailbox_1_s1,
                                  cpu_1_data_master_requests_mailbox_1_s1,
                                  cpu_2_data_master_granted_mailbox_1_s1,
                                  cpu_2_data_master_qualified_request_mailbox_1_s1,
                                  cpu_2_data_master_read_data_valid_mailbox_1_s1,
                                  cpu_2_data_master_requests_mailbox_1_s1,
                                  cpu_3_data_master_granted_mailbox_1_s1,
                                  cpu_3_data_master_qualified_request_mailbox_1_s1,
                                  cpu_3_data_master_read_data_valid_mailbox_1_s1,
                                  cpu_3_data_master_requests_mailbox_1_s1,
                                  d1_mailbox_1_s1_end_xfer,
                                  mailbox_1_s1_address,
                                  mailbox_1_s1_chipselect,
                                  mailbox_1_s1_read,
                                  mailbox_1_s1_readdata_from_sa,
                                  mailbox_1_s1_reset_n,
                                  mailbox_1_s1_write,
                                  mailbox_1_s1_writedata
                               )
;

  output           cpu_0_data_master_granted_mailbox_1_s1;
  output           cpu_0_data_master_qualified_request_mailbox_1_s1;
  output           cpu_0_data_master_read_data_valid_mailbox_1_s1;
  output           cpu_0_data_master_requests_mailbox_1_s1;
  output           cpu_1_data_master_granted_mailbox_1_s1;
  output           cpu_1_data_master_qualified_request_mailbox_1_s1;
  output           cpu_1_data_master_read_data_valid_mailbox_1_s1;
  output           cpu_1_data_master_requests_mailbox_1_s1;
  output           cpu_2_data_master_granted_mailbox_1_s1;
  output           cpu_2_data_master_qualified_request_mailbox_1_s1;
  output           cpu_2_data_master_read_data_valid_mailbox_1_s1;
  output           cpu_2_data_master_requests_mailbox_1_s1;
  output           cpu_3_data_master_granted_mailbox_1_s1;
  output           cpu_3_data_master_qualified_request_mailbox_1_s1;
  output           cpu_3_data_master_read_data_valid_mailbox_1_s1;
  output           cpu_3_data_master_requests_mailbox_1_s1;
  output           d1_mailbox_1_s1_end_xfer;
  output  [  1: 0] mailbox_1_s1_address;
  output           mailbox_1_s1_chipselect;
  output           mailbox_1_s1_read;
  output  [ 31: 0] mailbox_1_s1_readdata_from_sa;
  output           mailbox_1_s1_reset_n;
  output           mailbox_1_s1_write;
  output  [ 31: 0] mailbox_1_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 31: 0] mailbox_1_s1_readdata;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_mailbox_1_s1;
  wire             cpu_0_data_master_qualified_request_mailbox_1_s1;
  wire             cpu_0_data_master_read_data_valid_mailbox_1_s1;
  wire             cpu_0_data_master_requests_mailbox_1_s1;
  wire             cpu_0_data_master_saved_grant_mailbox_1_s1;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_mailbox_1_s1;
  wire             cpu_1_data_master_qualified_request_mailbox_1_s1;
  wire             cpu_1_data_master_read_data_valid_mailbox_1_s1;
  wire             cpu_1_data_master_requests_mailbox_1_s1;
  wire             cpu_1_data_master_saved_grant_mailbox_1_s1;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_mailbox_1_s1;
  wire             cpu_2_data_master_qualified_request_mailbox_1_s1;
  wire             cpu_2_data_master_read_data_valid_mailbox_1_s1;
  wire             cpu_2_data_master_requests_mailbox_1_s1;
  wire             cpu_2_data_master_saved_grant_mailbox_1_s1;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_mailbox_1_s1;
  wire             cpu_3_data_master_qualified_request_mailbox_1_s1;
  wire             cpu_3_data_master_read_data_valid_mailbox_1_s1;
  wire             cpu_3_data_master_requests_mailbox_1_s1;
  wire             cpu_3_data_master_saved_grant_mailbox_1_s1;
  reg              d1_mailbox_1_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_mailbox_1_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_mailbox_1_s1;
  reg              last_cycle_cpu_1_data_master_granted_slave_mailbox_1_s1;
  reg              last_cycle_cpu_2_data_master_granted_slave_mailbox_1_s1;
  reg              last_cycle_cpu_3_data_master_granted_slave_mailbox_1_s1;
  wire    [  1: 0] mailbox_1_s1_address;
  wire             mailbox_1_s1_allgrants;
  wire             mailbox_1_s1_allow_new_arb_cycle;
  wire             mailbox_1_s1_any_bursting_master_saved_grant;
  wire             mailbox_1_s1_any_continuerequest;
  reg     [  3: 0] mailbox_1_s1_arb_addend;
  wire             mailbox_1_s1_arb_counter_enable;
  reg     [  2: 0] mailbox_1_s1_arb_share_counter;
  wire    [  2: 0] mailbox_1_s1_arb_share_counter_next_value;
  wire    [  2: 0] mailbox_1_s1_arb_share_set_values;
  wire    [  3: 0] mailbox_1_s1_arb_winner;
  wire             mailbox_1_s1_arbitration_holdoff_internal;
  wire             mailbox_1_s1_beginbursttransfer_internal;
  wire             mailbox_1_s1_begins_xfer;
  wire             mailbox_1_s1_chipselect;
  wire    [  7: 0] mailbox_1_s1_chosen_master_double_vector;
  wire    [  3: 0] mailbox_1_s1_chosen_master_rot_left;
  wire             mailbox_1_s1_end_xfer;
  wire             mailbox_1_s1_firsttransfer;
  wire    [  3: 0] mailbox_1_s1_grant_vector;
  wire             mailbox_1_s1_in_a_read_cycle;
  wire             mailbox_1_s1_in_a_write_cycle;
  wire    [  3: 0] mailbox_1_s1_master_qreq_vector;
  wire             mailbox_1_s1_non_bursting_master_requests;
  wire             mailbox_1_s1_read;
  wire    [ 31: 0] mailbox_1_s1_readdata_from_sa;
  reg              mailbox_1_s1_reg_firsttransfer;
  wire             mailbox_1_s1_reset_n;
  reg     [  3: 0] mailbox_1_s1_saved_chosen_master_vector;
  reg              mailbox_1_s1_slavearbiterlockenable;
  wire             mailbox_1_s1_slavearbiterlockenable2;
  wire             mailbox_1_s1_unreg_firsttransfer;
  wire             mailbox_1_s1_waits_for_read;
  wire             mailbox_1_s1_waits_for_write;
  wire             mailbox_1_s1_write;
  wire    [ 31: 0] mailbox_1_s1_writedata;
  wire    [ 24: 0] shifted_address_to_mailbox_1_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_1_s1_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_1_s1_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_1_s1_from_cpu_3_data_master;
  wire             wait_for_mailbox_1_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~mailbox_1_s1_end_xfer;
    end


  assign mailbox_1_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_mailbox_1_s1 | cpu_1_data_master_qualified_request_mailbox_1_s1 | cpu_2_data_master_qualified_request_mailbox_1_s1 | cpu_3_data_master_qualified_request_mailbox_1_s1));
  //assign mailbox_1_s1_readdata_from_sa = mailbox_1_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign mailbox_1_s1_readdata_from_sa = mailbox_1_s1_readdata;

  assign cpu_0_data_master_requests_mailbox_1_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h50) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //mailbox_1_s1_arb_share_counter set values, which is an e_mux
  assign mailbox_1_s1_arb_share_set_values = 1;

  //mailbox_1_s1_non_bursting_master_requests mux, which is an e_mux
  assign mailbox_1_s1_non_bursting_master_requests = cpu_0_data_master_requests_mailbox_1_s1 |
    cpu_1_data_master_requests_mailbox_1_s1 |
    cpu_2_data_master_requests_mailbox_1_s1 |
    cpu_3_data_master_requests_mailbox_1_s1 |
    cpu_0_data_master_requests_mailbox_1_s1 |
    cpu_1_data_master_requests_mailbox_1_s1 |
    cpu_2_data_master_requests_mailbox_1_s1 |
    cpu_3_data_master_requests_mailbox_1_s1 |
    cpu_0_data_master_requests_mailbox_1_s1 |
    cpu_1_data_master_requests_mailbox_1_s1 |
    cpu_2_data_master_requests_mailbox_1_s1 |
    cpu_3_data_master_requests_mailbox_1_s1 |
    cpu_0_data_master_requests_mailbox_1_s1 |
    cpu_1_data_master_requests_mailbox_1_s1 |
    cpu_2_data_master_requests_mailbox_1_s1 |
    cpu_3_data_master_requests_mailbox_1_s1;

  //mailbox_1_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign mailbox_1_s1_any_bursting_master_saved_grant = 0;

  //mailbox_1_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign mailbox_1_s1_arb_share_counter_next_value = mailbox_1_s1_firsttransfer ? (mailbox_1_s1_arb_share_set_values - 1) : |mailbox_1_s1_arb_share_counter ? (mailbox_1_s1_arb_share_counter - 1) : 0;

  //mailbox_1_s1_allgrants all slave grants, which is an e_mux
  assign mailbox_1_s1_allgrants = (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector) |
    (|mailbox_1_s1_grant_vector);

  //mailbox_1_s1_end_xfer assignment, which is an e_assign
  assign mailbox_1_s1_end_xfer = ~(mailbox_1_s1_waits_for_read | mailbox_1_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_mailbox_1_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_mailbox_1_s1 = mailbox_1_s1_end_xfer & (~mailbox_1_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //mailbox_1_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign mailbox_1_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_mailbox_1_s1 & mailbox_1_s1_allgrants) | (end_xfer_arb_share_counter_term_mailbox_1_s1 & ~mailbox_1_s1_non_bursting_master_requests);

  //mailbox_1_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_1_s1_arb_share_counter <= 0;
      else if (mailbox_1_s1_arb_counter_enable)
          mailbox_1_s1_arb_share_counter <= mailbox_1_s1_arb_share_counter_next_value;
    end


  //mailbox_1_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_1_s1_slavearbiterlockenable <= 0;
      else if ((|mailbox_1_s1_master_qreq_vector & end_xfer_arb_share_counter_term_mailbox_1_s1) | (end_xfer_arb_share_counter_term_mailbox_1_s1 & ~mailbox_1_s1_non_bursting_master_requests))
          mailbox_1_s1_slavearbiterlockenable <= |mailbox_1_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master mailbox_1/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = mailbox_1_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //mailbox_1_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign mailbox_1_s1_slavearbiterlockenable2 = |mailbox_1_s1_arb_share_counter_next_value;

  //cpu_0/data_master mailbox_1/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = mailbox_1_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_1/data_master mailbox_1/s1 arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = mailbox_1_s1_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master mailbox_1/s1 arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = mailbox_1_s1_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted mailbox_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_mailbox_1_s1 <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_mailbox_1_s1 <= cpu_1_data_master_saved_grant_mailbox_1_s1 ? 1 : (mailbox_1_s1_arbitration_holdoff_internal | ~cpu_1_data_master_requests_mailbox_1_s1) ? 0 : last_cycle_cpu_1_data_master_granted_slave_mailbox_1_s1;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_mailbox_1_s1 & cpu_1_data_master_requests_mailbox_1_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_mailbox_1_s1 & cpu_1_data_master_requests_mailbox_1_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_mailbox_1_s1 & cpu_1_data_master_requests_mailbox_1_s1);

  //mailbox_1_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign mailbox_1_s1_any_continuerequest = cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest;

  //cpu_2/data_master mailbox_1/s1 arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = mailbox_1_s1_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master mailbox_1/s1 arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = mailbox_1_s1_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted mailbox_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_mailbox_1_s1 <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_mailbox_1_s1 <= cpu_2_data_master_saved_grant_mailbox_1_s1 ? 1 : (mailbox_1_s1_arbitration_holdoff_internal | ~cpu_2_data_master_requests_mailbox_1_s1) ? 0 : last_cycle_cpu_2_data_master_granted_slave_mailbox_1_s1;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_mailbox_1_s1 & cpu_2_data_master_requests_mailbox_1_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_mailbox_1_s1 & cpu_2_data_master_requests_mailbox_1_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_mailbox_1_s1 & cpu_2_data_master_requests_mailbox_1_s1);

  //cpu_3/data_master mailbox_1/s1 arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = mailbox_1_s1_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master mailbox_1/s1 arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = mailbox_1_s1_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted mailbox_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_mailbox_1_s1 <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_mailbox_1_s1 <= cpu_3_data_master_saved_grant_mailbox_1_s1 ? 1 : (mailbox_1_s1_arbitration_holdoff_internal | ~cpu_3_data_master_requests_mailbox_1_s1) ? 0 : last_cycle_cpu_3_data_master_granted_slave_mailbox_1_s1;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_mailbox_1_s1 & cpu_3_data_master_requests_mailbox_1_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_mailbox_1_s1 & cpu_3_data_master_requests_mailbox_1_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_mailbox_1_s1 & cpu_3_data_master_requests_mailbox_1_s1);

  assign cpu_0_data_master_qualified_request_mailbox_1_s1 = cpu_0_data_master_requests_mailbox_1_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_mailbox_1_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_mailbox_1_s1 = cpu_0_data_master_granted_mailbox_1_s1 & cpu_0_data_master_read & ~mailbox_1_s1_waits_for_read;

  //mailbox_1_s1_writedata mux, which is an e_mux
  assign mailbox_1_s1_writedata = (cpu_0_data_master_granted_mailbox_1_s1)? cpu_0_data_master_writedata :
    (cpu_1_data_master_granted_mailbox_1_s1)? cpu_1_data_master_writedata :
    (cpu_2_data_master_granted_mailbox_1_s1)? cpu_2_data_master_writedata :
    cpu_3_data_master_writedata;

  assign cpu_1_data_master_requests_mailbox_1_s1 = ({cpu_1_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h50) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //cpu_0/data_master granted mailbox_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_mailbox_1_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_mailbox_1_s1 <= cpu_0_data_master_saved_grant_mailbox_1_s1 ? 1 : (mailbox_1_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_mailbox_1_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_mailbox_1_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_mailbox_1_s1 & cpu_0_data_master_requests_mailbox_1_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_mailbox_1_s1 & cpu_0_data_master_requests_mailbox_1_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_mailbox_1_s1 & cpu_0_data_master_requests_mailbox_1_s1);

  assign cpu_1_data_master_qualified_request_mailbox_1_s1 = cpu_1_data_master_requests_mailbox_1_s1 & ~((cpu_1_data_master_read & ((cpu_1_data_master_latency_counter != 0) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_1_data_master_read_data_valid_mailbox_1_s1, which is an e_mux
  assign cpu_1_data_master_read_data_valid_mailbox_1_s1 = cpu_1_data_master_granted_mailbox_1_s1 & cpu_1_data_master_read & ~mailbox_1_s1_waits_for_read;

  assign cpu_2_data_master_requests_mailbox_1_s1 = ({cpu_2_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h50) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_mailbox_1_s1 = cpu_2_data_master_requests_mailbox_1_s1 & ~((cpu_2_data_master_read & ((cpu_2_data_master_latency_counter != 0) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_2_data_master_read_data_valid_mailbox_1_s1, which is an e_mux
  assign cpu_2_data_master_read_data_valid_mailbox_1_s1 = cpu_2_data_master_granted_mailbox_1_s1 & cpu_2_data_master_read & ~mailbox_1_s1_waits_for_read;

  assign cpu_3_data_master_requests_mailbox_1_s1 = ({cpu_3_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h50) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_mailbox_1_s1 = cpu_3_data_master_requests_mailbox_1_s1 & ~((cpu_3_data_master_read & ((cpu_3_data_master_latency_counter != 0) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock);
  //local readdatavalid cpu_3_data_master_read_data_valid_mailbox_1_s1, which is an e_mux
  assign cpu_3_data_master_read_data_valid_mailbox_1_s1 = cpu_3_data_master_granted_mailbox_1_s1 & cpu_3_data_master_read & ~mailbox_1_s1_waits_for_read;

  //allow new arb cycle for mailbox_1/s1, which is an e_assign
  assign mailbox_1_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_3_data_master_arbiterlock;

  //cpu_3/data_master assignment into master qualified-requests vector for mailbox_1/s1, which is an e_assign
  assign mailbox_1_s1_master_qreq_vector[0] = cpu_3_data_master_qualified_request_mailbox_1_s1;

  //cpu_3/data_master grant mailbox_1/s1, which is an e_assign
  assign cpu_3_data_master_granted_mailbox_1_s1 = mailbox_1_s1_grant_vector[0];

  //cpu_3/data_master saved-grant mailbox_1/s1, which is an e_assign
  assign cpu_3_data_master_saved_grant_mailbox_1_s1 = mailbox_1_s1_arb_winner[0] && cpu_3_data_master_requests_mailbox_1_s1;

  //cpu_2/data_master assignment into master qualified-requests vector for mailbox_1/s1, which is an e_assign
  assign mailbox_1_s1_master_qreq_vector[1] = cpu_2_data_master_qualified_request_mailbox_1_s1;

  //cpu_2/data_master grant mailbox_1/s1, which is an e_assign
  assign cpu_2_data_master_granted_mailbox_1_s1 = mailbox_1_s1_grant_vector[1];

  //cpu_2/data_master saved-grant mailbox_1/s1, which is an e_assign
  assign cpu_2_data_master_saved_grant_mailbox_1_s1 = mailbox_1_s1_arb_winner[1] && cpu_2_data_master_requests_mailbox_1_s1;

  //cpu_1/data_master assignment into master qualified-requests vector for mailbox_1/s1, which is an e_assign
  assign mailbox_1_s1_master_qreq_vector[2] = cpu_1_data_master_qualified_request_mailbox_1_s1;

  //cpu_1/data_master grant mailbox_1/s1, which is an e_assign
  assign cpu_1_data_master_granted_mailbox_1_s1 = mailbox_1_s1_grant_vector[2];

  //cpu_1/data_master saved-grant mailbox_1/s1, which is an e_assign
  assign cpu_1_data_master_saved_grant_mailbox_1_s1 = mailbox_1_s1_arb_winner[2] && cpu_1_data_master_requests_mailbox_1_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for mailbox_1/s1, which is an e_assign
  assign mailbox_1_s1_master_qreq_vector[3] = cpu_0_data_master_qualified_request_mailbox_1_s1;

  //cpu_0/data_master grant mailbox_1/s1, which is an e_assign
  assign cpu_0_data_master_granted_mailbox_1_s1 = mailbox_1_s1_grant_vector[3];

  //cpu_0/data_master saved-grant mailbox_1/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_mailbox_1_s1 = mailbox_1_s1_arb_winner[3] && cpu_0_data_master_requests_mailbox_1_s1;

  //mailbox_1/s1 chosen-master double-vector, which is an e_assign
  assign mailbox_1_s1_chosen_master_double_vector = {mailbox_1_s1_master_qreq_vector, mailbox_1_s1_master_qreq_vector} & ({~mailbox_1_s1_master_qreq_vector, ~mailbox_1_s1_master_qreq_vector} + mailbox_1_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign mailbox_1_s1_arb_winner = (mailbox_1_s1_allow_new_arb_cycle & | mailbox_1_s1_grant_vector) ? mailbox_1_s1_grant_vector : mailbox_1_s1_saved_chosen_master_vector;

  //saved mailbox_1_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_1_s1_saved_chosen_master_vector <= 0;
      else if (mailbox_1_s1_allow_new_arb_cycle)
          mailbox_1_s1_saved_chosen_master_vector <= |mailbox_1_s1_grant_vector ? mailbox_1_s1_grant_vector : mailbox_1_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign mailbox_1_s1_grant_vector = {(mailbox_1_s1_chosen_master_double_vector[3] | mailbox_1_s1_chosen_master_double_vector[7]),
    (mailbox_1_s1_chosen_master_double_vector[2] | mailbox_1_s1_chosen_master_double_vector[6]),
    (mailbox_1_s1_chosen_master_double_vector[1] | mailbox_1_s1_chosen_master_double_vector[5]),
    (mailbox_1_s1_chosen_master_double_vector[0] | mailbox_1_s1_chosen_master_double_vector[4])};

  //mailbox_1/s1 chosen master rotated left, which is an e_assign
  assign mailbox_1_s1_chosen_master_rot_left = (mailbox_1_s1_arb_winner << 1) ? (mailbox_1_s1_arb_winner << 1) : 1;

  //mailbox_1/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_1_s1_arb_addend <= 1;
      else if (|mailbox_1_s1_grant_vector)
          mailbox_1_s1_arb_addend <= mailbox_1_s1_end_xfer? mailbox_1_s1_chosen_master_rot_left : mailbox_1_s1_grant_vector;
    end


  //mailbox_1_s1_reset_n assignment, which is an e_assign
  assign mailbox_1_s1_reset_n = reset_n;

  assign mailbox_1_s1_chipselect = cpu_0_data_master_granted_mailbox_1_s1 | cpu_1_data_master_granted_mailbox_1_s1 | cpu_2_data_master_granted_mailbox_1_s1 | cpu_3_data_master_granted_mailbox_1_s1;
  //mailbox_1_s1_firsttransfer first transaction, which is an e_assign
  assign mailbox_1_s1_firsttransfer = mailbox_1_s1_begins_xfer ? mailbox_1_s1_unreg_firsttransfer : mailbox_1_s1_reg_firsttransfer;

  //mailbox_1_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign mailbox_1_s1_unreg_firsttransfer = ~(mailbox_1_s1_slavearbiterlockenable & mailbox_1_s1_any_continuerequest);

  //mailbox_1_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_1_s1_reg_firsttransfer <= 1'b1;
      else if (mailbox_1_s1_begins_xfer)
          mailbox_1_s1_reg_firsttransfer <= mailbox_1_s1_unreg_firsttransfer;
    end


  //mailbox_1_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign mailbox_1_s1_beginbursttransfer_internal = mailbox_1_s1_begins_xfer;

  //mailbox_1_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign mailbox_1_s1_arbitration_holdoff_internal = mailbox_1_s1_begins_xfer & mailbox_1_s1_firsttransfer;

  //mailbox_1_s1_read assignment, which is an e_mux
  assign mailbox_1_s1_read = (cpu_0_data_master_granted_mailbox_1_s1 & cpu_0_data_master_read) | (cpu_1_data_master_granted_mailbox_1_s1 & cpu_1_data_master_read) | (cpu_2_data_master_granted_mailbox_1_s1 & cpu_2_data_master_read) | (cpu_3_data_master_granted_mailbox_1_s1 & cpu_3_data_master_read);

  //mailbox_1_s1_write assignment, which is an e_mux
  assign mailbox_1_s1_write = (cpu_0_data_master_granted_mailbox_1_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_mailbox_1_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_mailbox_1_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_mailbox_1_s1 & cpu_3_data_master_write);

  assign shifted_address_to_mailbox_1_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //mailbox_1_s1_address mux, which is an e_mux
  assign mailbox_1_s1_address = (cpu_0_data_master_granted_mailbox_1_s1)? (shifted_address_to_mailbox_1_s1_from_cpu_0_data_master >> 2) :
    (cpu_1_data_master_granted_mailbox_1_s1)? (shifted_address_to_mailbox_1_s1_from_cpu_1_data_master >> 2) :
    (cpu_2_data_master_granted_mailbox_1_s1)? (shifted_address_to_mailbox_1_s1_from_cpu_2_data_master >> 2) :
    (shifted_address_to_mailbox_1_s1_from_cpu_3_data_master >> 2);

  assign shifted_address_to_mailbox_1_s1_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_mailbox_1_s1_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_mailbox_1_s1_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  //d1_mailbox_1_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_mailbox_1_s1_end_xfer <= 1;
      else 
        d1_mailbox_1_s1_end_xfer <= mailbox_1_s1_end_xfer;
    end


  //mailbox_1_s1_waits_for_read in a cycle, which is an e_mux
  assign mailbox_1_s1_waits_for_read = mailbox_1_s1_in_a_read_cycle & mailbox_1_s1_begins_xfer;

  //mailbox_1_s1_in_a_read_cycle assignment, which is an e_assign
  assign mailbox_1_s1_in_a_read_cycle = (cpu_0_data_master_granted_mailbox_1_s1 & cpu_0_data_master_read) | (cpu_1_data_master_granted_mailbox_1_s1 & cpu_1_data_master_read) | (cpu_2_data_master_granted_mailbox_1_s1 & cpu_2_data_master_read) | (cpu_3_data_master_granted_mailbox_1_s1 & cpu_3_data_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = mailbox_1_s1_in_a_read_cycle;

  //mailbox_1_s1_waits_for_write in a cycle, which is an e_mux
  assign mailbox_1_s1_waits_for_write = mailbox_1_s1_in_a_write_cycle & 0;

  //mailbox_1_s1_in_a_write_cycle assignment, which is an e_assign
  assign mailbox_1_s1_in_a_write_cycle = (cpu_0_data_master_granted_mailbox_1_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_mailbox_1_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_mailbox_1_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_mailbox_1_s1 & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = mailbox_1_s1_in_a_write_cycle;

  assign wait_for_mailbox_1_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //mailbox_1/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_mailbox_1_s1 + cpu_1_data_master_granted_mailbox_1_s1 + cpu_2_data_master_granted_mailbox_1_s1 + cpu_3_data_master_granted_mailbox_1_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_mailbox_1_s1 + cpu_1_data_master_saved_grant_mailbox_1_s1 + cpu_2_data_master_saved_grant_mailbox_1_s1 + cpu_3_data_master_saved_grant_mailbox_1_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module mailbox_2_s1_arbitrator (
                                 // inputs:
                                  clk,
                                  cpu_0_data_master_address_to_slave,
                                  cpu_0_data_master_latency_counter,
                                  cpu_0_data_master_read,
                                  cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_0_data_master_write,
                                  cpu_0_data_master_writedata,
                                  cpu_1_data_master_address_to_slave,
                                  cpu_1_data_master_latency_counter,
                                  cpu_1_data_master_read,
                                  cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_1_data_master_write,
                                  cpu_1_data_master_writedata,
                                  cpu_2_data_master_address_to_slave,
                                  cpu_2_data_master_latency_counter,
                                  cpu_2_data_master_read,
                                  cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_2_data_master_write,
                                  cpu_2_data_master_writedata,
                                  cpu_3_data_master_address_to_slave,
                                  cpu_3_data_master_latency_counter,
                                  cpu_3_data_master_read,
                                  cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_3_data_master_write,
                                  cpu_3_data_master_writedata,
                                  mailbox_2_s1_readdata,
                                  reset_n,

                                 // outputs:
                                  cpu_0_data_master_granted_mailbox_2_s1,
                                  cpu_0_data_master_qualified_request_mailbox_2_s1,
                                  cpu_0_data_master_read_data_valid_mailbox_2_s1,
                                  cpu_0_data_master_requests_mailbox_2_s1,
                                  cpu_1_data_master_granted_mailbox_2_s1,
                                  cpu_1_data_master_qualified_request_mailbox_2_s1,
                                  cpu_1_data_master_read_data_valid_mailbox_2_s1,
                                  cpu_1_data_master_requests_mailbox_2_s1,
                                  cpu_2_data_master_granted_mailbox_2_s1,
                                  cpu_2_data_master_qualified_request_mailbox_2_s1,
                                  cpu_2_data_master_read_data_valid_mailbox_2_s1,
                                  cpu_2_data_master_requests_mailbox_2_s1,
                                  cpu_3_data_master_granted_mailbox_2_s1,
                                  cpu_3_data_master_qualified_request_mailbox_2_s1,
                                  cpu_3_data_master_read_data_valid_mailbox_2_s1,
                                  cpu_3_data_master_requests_mailbox_2_s1,
                                  d1_mailbox_2_s1_end_xfer,
                                  mailbox_2_s1_address,
                                  mailbox_2_s1_chipselect,
                                  mailbox_2_s1_read,
                                  mailbox_2_s1_readdata_from_sa,
                                  mailbox_2_s1_reset_n,
                                  mailbox_2_s1_write,
                                  mailbox_2_s1_writedata
                               )
;

  output           cpu_0_data_master_granted_mailbox_2_s1;
  output           cpu_0_data_master_qualified_request_mailbox_2_s1;
  output           cpu_0_data_master_read_data_valid_mailbox_2_s1;
  output           cpu_0_data_master_requests_mailbox_2_s1;
  output           cpu_1_data_master_granted_mailbox_2_s1;
  output           cpu_1_data_master_qualified_request_mailbox_2_s1;
  output           cpu_1_data_master_read_data_valid_mailbox_2_s1;
  output           cpu_1_data_master_requests_mailbox_2_s1;
  output           cpu_2_data_master_granted_mailbox_2_s1;
  output           cpu_2_data_master_qualified_request_mailbox_2_s1;
  output           cpu_2_data_master_read_data_valid_mailbox_2_s1;
  output           cpu_2_data_master_requests_mailbox_2_s1;
  output           cpu_3_data_master_granted_mailbox_2_s1;
  output           cpu_3_data_master_qualified_request_mailbox_2_s1;
  output           cpu_3_data_master_read_data_valid_mailbox_2_s1;
  output           cpu_3_data_master_requests_mailbox_2_s1;
  output           d1_mailbox_2_s1_end_xfer;
  output  [  1: 0] mailbox_2_s1_address;
  output           mailbox_2_s1_chipselect;
  output           mailbox_2_s1_read;
  output  [ 31: 0] mailbox_2_s1_readdata_from_sa;
  output           mailbox_2_s1_reset_n;
  output           mailbox_2_s1_write;
  output  [ 31: 0] mailbox_2_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 31: 0] mailbox_2_s1_readdata;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_mailbox_2_s1;
  wire             cpu_0_data_master_qualified_request_mailbox_2_s1;
  wire             cpu_0_data_master_read_data_valid_mailbox_2_s1;
  wire             cpu_0_data_master_requests_mailbox_2_s1;
  wire             cpu_0_data_master_saved_grant_mailbox_2_s1;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_mailbox_2_s1;
  wire             cpu_1_data_master_qualified_request_mailbox_2_s1;
  wire             cpu_1_data_master_read_data_valid_mailbox_2_s1;
  wire             cpu_1_data_master_requests_mailbox_2_s1;
  wire             cpu_1_data_master_saved_grant_mailbox_2_s1;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_mailbox_2_s1;
  wire             cpu_2_data_master_qualified_request_mailbox_2_s1;
  wire             cpu_2_data_master_read_data_valid_mailbox_2_s1;
  wire             cpu_2_data_master_requests_mailbox_2_s1;
  wire             cpu_2_data_master_saved_grant_mailbox_2_s1;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_mailbox_2_s1;
  wire             cpu_3_data_master_qualified_request_mailbox_2_s1;
  wire             cpu_3_data_master_read_data_valid_mailbox_2_s1;
  wire             cpu_3_data_master_requests_mailbox_2_s1;
  wire             cpu_3_data_master_saved_grant_mailbox_2_s1;
  reg              d1_mailbox_2_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_mailbox_2_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_mailbox_2_s1;
  reg              last_cycle_cpu_1_data_master_granted_slave_mailbox_2_s1;
  reg              last_cycle_cpu_2_data_master_granted_slave_mailbox_2_s1;
  reg              last_cycle_cpu_3_data_master_granted_slave_mailbox_2_s1;
  wire    [  1: 0] mailbox_2_s1_address;
  wire             mailbox_2_s1_allgrants;
  wire             mailbox_2_s1_allow_new_arb_cycle;
  wire             mailbox_2_s1_any_bursting_master_saved_grant;
  wire             mailbox_2_s1_any_continuerequest;
  reg     [  3: 0] mailbox_2_s1_arb_addend;
  wire             mailbox_2_s1_arb_counter_enable;
  reg     [  2: 0] mailbox_2_s1_arb_share_counter;
  wire    [  2: 0] mailbox_2_s1_arb_share_counter_next_value;
  wire    [  2: 0] mailbox_2_s1_arb_share_set_values;
  wire    [  3: 0] mailbox_2_s1_arb_winner;
  wire             mailbox_2_s1_arbitration_holdoff_internal;
  wire             mailbox_2_s1_beginbursttransfer_internal;
  wire             mailbox_2_s1_begins_xfer;
  wire             mailbox_2_s1_chipselect;
  wire    [  7: 0] mailbox_2_s1_chosen_master_double_vector;
  wire    [  3: 0] mailbox_2_s1_chosen_master_rot_left;
  wire             mailbox_2_s1_end_xfer;
  wire             mailbox_2_s1_firsttransfer;
  wire    [  3: 0] mailbox_2_s1_grant_vector;
  wire             mailbox_2_s1_in_a_read_cycle;
  wire             mailbox_2_s1_in_a_write_cycle;
  wire    [  3: 0] mailbox_2_s1_master_qreq_vector;
  wire             mailbox_2_s1_non_bursting_master_requests;
  wire             mailbox_2_s1_read;
  wire    [ 31: 0] mailbox_2_s1_readdata_from_sa;
  reg              mailbox_2_s1_reg_firsttransfer;
  wire             mailbox_2_s1_reset_n;
  reg     [  3: 0] mailbox_2_s1_saved_chosen_master_vector;
  reg              mailbox_2_s1_slavearbiterlockenable;
  wire             mailbox_2_s1_slavearbiterlockenable2;
  wire             mailbox_2_s1_unreg_firsttransfer;
  wire             mailbox_2_s1_waits_for_read;
  wire             mailbox_2_s1_waits_for_write;
  wire             mailbox_2_s1_write;
  wire    [ 31: 0] mailbox_2_s1_writedata;
  wire    [ 24: 0] shifted_address_to_mailbox_2_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_2_s1_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_2_s1_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_2_s1_from_cpu_3_data_master;
  wire             wait_for_mailbox_2_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~mailbox_2_s1_end_xfer;
    end


  assign mailbox_2_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_mailbox_2_s1 | cpu_1_data_master_qualified_request_mailbox_2_s1 | cpu_2_data_master_qualified_request_mailbox_2_s1 | cpu_3_data_master_qualified_request_mailbox_2_s1));
  //assign mailbox_2_s1_readdata_from_sa = mailbox_2_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign mailbox_2_s1_readdata_from_sa = mailbox_2_s1_readdata;

  assign cpu_0_data_master_requests_mailbox_2_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h70) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //mailbox_2_s1_arb_share_counter set values, which is an e_mux
  assign mailbox_2_s1_arb_share_set_values = 1;

  //mailbox_2_s1_non_bursting_master_requests mux, which is an e_mux
  assign mailbox_2_s1_non_bursting_master_requests = cpu_0_data_master_requests_mailbox_2_s1 |
    cpu_1_data_master_requests_mailbox_2_s1 |
    cpu_2_data_master_requests_mailbox_2_s1 |
    cpu_3_data_master_requests_mailbox_2_s1 |
    cpu_0_data_master_requests_mailbox_2_s1 |
    cpu_1_data_master_requests_mailbox_2_s1 |
    cpu_2_data_master_requests_mailbox_2_s1 |
    cpu_3_data_master_requests_mailbox_2_s1 |
    cpu_0_data_master_requests_mailbox_2_s1 |
    cpu_1_data_master_requests_mailbox_2_s1 |
    cpu_2_data_master_requests_mailbox_2_s1 |
    cpu_3_data_master_requests_mailbox_2_s1 |
    cpu_0_data_master_requests_mailbox_2_s1 |
    cpu_1_data_master_requests_mailbox_2_s1 |
    cpu_2_data_master_requests_mailbox_2_s1 |
    cpu_3_data_master_requests_mailbox_2_s1;

  //mailbox_2_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign mailbox_2_s1_any_bursting_master_saved_grant = 0;

  //mailbox_2_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign mailbox_2_s1_arb_share_counter_next_value = mailbox_2_s1_firsttransfer ? (mailbox_2_s1_arb_share_set_values - 1) : |mailbox_2_s1_arb_share_counter ? (mailbox_2_s1_arb_share_counter - 1) : 0;

  //mailbox_2_s1_allgrants all slave grants, which is an e_mux
  assign mailbox_2_s1_allgrants = (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector) |
    (|mailbox_2_s1_grant_vector);

  //mailbox_2_s1_end_xfer assignment, which is an e_assign
  assign mailbox_2_s1_end_xfer = ~(mailbox_2_s1_waits_for_read | mailbox_2_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_mailbox_2_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_mailbox_2_s1 = mailbox_2_s1_end_xfer & (~mailbox_2_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //mailbox_2_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign mailbox_2_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_mailbox_2_s1 & mailbox_2_s1_allgrants) | (end_xfer_arb_share_counter_term_mailbox_2_s1 & ~mailbox_2_s1_non_bursting_master_requests);

  //mailbox_2_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_2_s1_arb_share_counter <= 0;
      else if (mailbox_2_s1_arb_counter_enable)
          mailbox_2_s1_arb_share_counter <= mailbox_2_s1_arb_share_counter_next_value;
    end


  //mailbox_2_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_2_s1_slavearbiterlockenable <= 0;
      else if ((|mailbox_2_s1_master_qreq_vector & end_xfer_arb_share_counter_term_mailbox_2_s1) | (end_xfer_arb_share_counter_term_mailbox_2_s1 & ~mailbox_2_s1_non_bursting_master_requests))
          mailbox_2_s1_slavearbiterlockenable <= |mailbox_2_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master mailbox_2/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = mailbox_2_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //mailbox_2_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign mailbox_2_s1_slavearbiterlockenable2 = |mailbox_2_s1_arb_share_counter_next_value;

  //cpu_0/data_master mailbox_2/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = mailbox_2_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_1/data_master mailbox_2/s1 arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = mailbox_2_s1_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master mailbox_2/s1 arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = mailbox_2_s1_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted mailbox_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_mailbox_2_s1 <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_mailbox_2_s1 <= cpu_1_data_master_saved_grant_mailbox_2_s1 ? 1 : (mailbox_2_s1_arbitration_holdoff_internal | ~cpu_1_data_master_requests_mailbox_2_s1) ? 0 : last_cycle_cpu_1_data_master_granted_slave_mailbox_2_s1;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_mailbox_2_s1 & cpu_1_data_master_requests_mailbox_2_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_mailbox_2_s1 & cpu_1_data_master_requests_mailbox_2_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_mailbox_2_s1 & cpu_1_data_master_requests_mailbox_2_s1);

  //mailbox_2_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign mailbox_2_s1_any_continuerequest = cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest;

  //cpu_2/data_master mailbox_2/s1 arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = mailbox_2_s1_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master mailbox_2/s1 arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = mailbox_2_s1_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted mailbox_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_mailbox_2_s1 <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_mailbox_2_s1 <= cpu_2_data_master_saved_grant_mailbox_2_s1 ? 1 : (mailbox_2_s1_arbitration_holdoff_internal | ~cpu_2_data_master_requests_mailbox_2_s1) ? 0 : last_cycle_cpu_2_data_master_granted_slave_mailbox_2_s1;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_mailbox_2_s1 & cpu_2_data_master_requests_mailbox_2_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_mailbox_2_s1 & cpu_2_data_master_requests_mailbox_2_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_mailbox_2_s1 & cpu_2_data_master_requests_mailbox_2_s1);

  //cpu_3/data_master mailbox_2/s1 arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = mailbox_2_s1_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master mailbox_2/s1 arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = mailbox_2_s1_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted mailbox_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_mailbox_2_s1 <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_mailbox_2_s1 <= cpu_3_data_master_saved_grant_mailbox_2_s1 ? 1 : (mailbox_2_s1_arbitration_holdoff_internal | ~cpu_3_data_master_requests_mailbox_2_s1) ? 0 : last_cycle_cpu_3_data_master_granted_slave_mailbox_2_s1;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_mailbox_2_s1 & cpu_3_data_master_requests_mailbox_2_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_mailbox_2_s1 & cpu_3_data_master_requests_mailbox_2_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_mailbox_2_s1 & cpu_3_data_master_requests_mailbox_2_s1);

  assign cpu_0_data_master_qualified_request_mailbox_2_s1 = cpu_0_data_master_requests_mailbox_2_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_mailbox_2_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_mailbox_2_s1 = cpu_0_data_master_granted_mailbox_2_s1 & cpu_0_data_master_read & ~mailbox_2_s1_waits_for_read;

  //mailbox_2_s1_writedata mux, which is an e_mux
  assign mailbox_2_s1_writedata = (cpu_0_data_master_granted_mailbox_2_s1)? cpu_0_data_master_writedata :
    (cpu_1_data_master_granted_mailbox_2_s1)? cpu_1_data_master_writedata :
    (cpu_2_data_master_granted_mailbox_2_s1)? cpu_2_data_master_writedata :
    cpu_3_data_master_writedata;

  assign cpu_1_data_master_requests_mailbox_2_s1 = ({cpu_1_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h70) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //cpu_0/data_master granted mailbox_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_mailbox_2_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_mailbox_2_s1 <= cpu_0_data_master_saved_grant_mailbox_2_s1 ? 1 : (mailbox_2_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_mailbox_2_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_mailbox_2_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_mailbox_2_s1 & cpu_0_data_master_requests_mailbox_2_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_mailbox_2_s1 & cpu_0_data_master_requests_mailbox_2_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_mailbox_2_s1 & cpu_0_data_master_requests_mailbox_2_s1);

  assign cpu_1_data_master_qualified_request_mailbox_2_s1 = cpu_1_data_master_requests_mailbox_2_s1 & ~((cpu_1_data_master_read & ((cpu_1_data_master_latency_counter != 0) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_1_data_master_read_data_valid_mailbox_2_s1, which is an e_mux
  assign cpu_1_data_master_read_data_valid_mailbox_2_s1 = cpu_1_data_master_granted_mailbox_2_s1 & cpu_1_data_master_read & ~mailbox_2_s1_waits_for_read;

  assign cpu_2_data_master_requests_mailbox_2_s1 = ({cpu_2_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h70) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_mailbox_2_s1 = cpu_2_data_master_requests_mailbox_2_s1 & ~((cpu_2_data_master_read & ((cpu_2_data_master_latency_counter != 0) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_2_data_master_read_data_valid_mailbox_2_s1, which is an e_mux
  assign cpu_2_data_master_read_data_valid_mailbox_2_s1 = cpu_2_data_master_granted_mailbox_2_s1 & cpu_2_data_master_read & ~mailbox_2_s1_waits_for_read;

  assign cpu_3_data_master_requests_mailbox_2_s1 = ({cpu_3_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h70) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_mailbox_2_s1 = cpu_3_data_master_requests_mailbox_2_s1 & ~((cpu_3_data_master_read & ((cpu_3_data_master_latency_counter != 0) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock);
  //local readdatavalid cpu_3_data_master_read_data_valid_mailbox_2_s1, which is an e_mux
  assign cpu_3_data_master_read_data_valid_mailbox_2_s1 = cpu_3_data_master_granted_mailbox_2_s1 & cpu_3_data_master_read & ~mailbox_2_s1_waits_for_read;

  //allow new arb cycle for mailbox_2/s1, which is an e_assign
  assign mailbox_2_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_3_data_master_arbiterlock;

  //cpu_3/data_master assignment into master qualified-requests vector for mailbox_2/s1, which is an e_assign
  assign mailbox_2_s1_master_qreq_vector[0] = cpu_3_data_master_qualified_request_mailbox_2_s1;

  //cpu_3/data_master grant mailbox_2/s1, which is an e_assign
  assign cpu_3_data_master_granted_mailbox_2_s1 = mailbox_2_s1_grant_vector[0];

  //cpu_3/data_master saved-grant mailbox_2/s1, which is an e_assign
  assign cpu_3_data_master_saved_grant_mailbox_2_s1 = mailbox_2_s1_arb_winner[0] && cpu_3_data_master_requests_mailbox_2_s1;

  //cpu_2/data_master assignment into master qualified-requests vector for mailbox_2/s1, which is an e_assign
  assign mailbox_2_s1_master_qreq_vector[1] = cpu_2_data_master_qualified_request_mailbox_2_s1;

  //cpu_2/data_master grant mailbox_2/s1, which is an e_assign
  assign cpu_2_data_master_granted_mailbox_2_s1 = mailbox_2_s1_grant_vector[1];

  //cpu_2/data_master saved-grant mailbox_2/s1, which is an e_assign
  assign cpu_2_data_master_saved_grant_mailbox_2_s1 = mailbox_2_s1_arb_winner[1] && cpu_2_data_master_requests_mailbox_2_s1;

  //cpu_1/data_master assignment into master qualified-requests vector for mailbox_2/s1, which is an e_assign
  assign mailbox_2_s1_master_qreq_vector[2] = cpu_1_data_master_qualified_request_mailbox_2_s1;

  //cpu_1/data_master grant mailbox_2/s1, which is an e_assign
  assign cpu_1_data_master_granted_mailbox_2_s1 = mailbox_2_s1_grant_vector[2];

  //cpu_1/data_master saved-grant mailbox_2/s1, which is an e_assign
  assign cpu_1_data_master_saved_grant_mailbox_2_s1 = mailbox_2_s1_arb_winner[2] && cpu_1_data_master_requests_mailbox_2_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for mailbox_2/s1, which is an e_assign
  assign mailbox_2_s1_master_qreq_vector[3] = cpu_0_data_master_qualified_request_mailbox_2_s1;

  //cpu_0/data_master grant mailbox_2/s1, which is an e_assign
  assign cpu_0_data_master_granted_mailbox_2_s1 = mailbox_2_s1_grant_vector[3];

  //cpu_0/data_master saved-grant mailbox_2/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_mailbox_2_s1 = mailbox_2_s1_arb_winner[3] && cpu_0_data_master_requests_mailbox_2_s1;

  //mailbox_2/s1 chosen-master double-vector, which is an e_assign
  assign mailbox_2_s1_chosen_master_double_vector = {mailbox_2_s1_master_qreq_vector, mailbox_2_s1_master_qreq_vector} & ({~mailbox_2_s1_master_qreq_vector, ~mailbox_2_s1_master_qreq_vector} + mailbox_2_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign mailbox_2_s1_arb_winner = (mailbox_2_s1_allow_new_arb_cycle & | mailbox_2_s1_grant_vector) ? mailbox_2_s1_grant_vector : mailbox_2_s1_saved_chosen_master_vector;

  //saved mailbox_2_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_2_s1_saved_chosen_master_vector <= 0;
      else if (mailbox_2_s1_allow_new_arb_cycle)
          mailbox_2_s1_saved_chosen_master_vector <= |mailbox_2_s1_grant_vector ? mailbox_2_s1_grant_vector : mailbox_2_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign mailbox_2_s1_grant_vector = {(mailbox_2_s1_chosen_master_double_vector[3] | mailbox_2_s1_chosen_master_double_vector[7]),
    (mailbox_2_s1_chosen_master_double_vector[2] | mailbox_2_s1_chosen_master_double_vector[6]),
    (mailbox_2_s1_chosen_master_double_vector[1] | mailbox_2_s1_chosen_master_double_vector[5]),
    (mailbox_2_s1_chosen_master_double_vector[0] | mailbox_2_s1_chosen_master_double_vector[4])};

  //mailbox_2/s1 chosen master rotated left, which is an e_assign
  assign mailbox_2_s1_chosen_master_rot_left = (mailbox_2_s1_arb_winner << 1) ? (mailbox_2_s1_arb_winner << 1) : 1;

  //mailbox_2/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_2_s1_arb_addend <= 1;
      else if (|mailbox_2_s1_grant_vector)
          mailbox_2_s1_arb_addend <= mailbox_2_s1_end_xfer? mailbox_2_s1_chosen_master_rot_left : mailbox_2_s1_grant_vector;
    end


  //mailbox_2_s1_reset_n assignment, which is an e_assign
  assign mailbox_2_s1_reset_n = reset_n;

  assign mailbox_2_s1_chipselect = cpu_0_data_master_granted_mailbox_2_s1 | cpu_1_data_master_granted_mailbox_2_s1 | cpu_2_data_master_granted_mailbox_2_s1 | cpu_3_data_master_granted_mailbox_2_s1;
  //mailbox_2_s1_firsttransfer first transaction, which is an e_assign
  assign mailbox_2_s1_firsttransfer = mailbox_2_s1_begins_xfer ? mailbox_2_s1_unreg_firsttransfer : mailbox_2_s1_reg_firsttransfer;

  //mailbox_2_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign mailbox_2_s1_unreg_firsttransfer = ~(mailbox_2_s1_slavearbiterlockenable & mailbox_2_s1_any_continuerequest);

  //mailbox_2_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_2_s1_reg_firsttransfer <= 1'b1;
      else if (mailbox_2_s1_begins_xfer)
          mailbox_2_s1_reg_firsttransfer <= mailbox_2_s1_unreg_firsttransfer;
    end


  //mailbox_2_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign mailbox_2_s1_beginbursttransfer_internal = mailbox_2_s1_begins_xfer;

  //mailbox_2_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign mailbox_2_s1_arbitration_holdoff_internal = mailbox_2_s1_begins_xfer & mailbox_2_s1_firsttransfer;

  //mailbox_2_s1_read assignment, which is an e_mux
  assign mailbox_2_s1_read = (cpu_0_data_master_granted_mailbox_2_s1 & cpu_0_data_master_read) | (cpu_1_data_master_granted_mailbox_2_s1 & cpu_1_data_master_read) | (cpu_2_data_master_granted_mailbox_2_s1 & cpu_2_data_master_read) | (cpu_3_data_master_granted_mailbox_2_s1 & cpu_3_data_master_read);

  //mailbox_2_s1_write assignment, which is an e_mux
  assign mailbox_2_s1_write = (cpu_0_data_master_granted_mailbox_2_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_mailbox_2_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_mailbox_2_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_mailbox_2_s1 & cpu_3_data_master_write);

  assign shifted_address_to_mailbox_2_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //mailbox_2_s1_address mux, which is an e_mux
  assign mailbox_2_s1_address = (cpu_0_data_master_granted_mailbox_2_s1)? (shifted_address_to_mailbox_2_s1_from_cpu_0_data_master >> 2) :
    (cpu_1_data_master_granted_mailbox_2_s1)? (shifted_address_to_mailbox_2_s1_from_cpu_1_data_master >> 2) :
    (cpu_2_data_master_granted_mailbox_2_s1)? (shifted_address_to_mailbox_2_s1_from_cpu_2_data_master >> 2) :
    (shifted_address_to_mailbox_2_s1_from_cpu_3_data_master >> 2);

  assign shifted_address_to_mailbox_2_s1_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_mailbox_2_s1_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_mailbox_2_s1_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  //d1_mailbox_2_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_mailbox_2_s1_end_xfer <= 1;
      else 
        d1_mailbox_2_s1_end_xfer <= mailbox_2_s1_end_xfer;
    end


  //mailbox_2_s1_waits_for_read in a cycle, which is an e_mux
  assign mailbox_2_s1_waits_for_read = mailbox_2_s1_in_a_read_cycle & mailbox_2_s1_begins_xfer;

  //mailbox_2_s1_in_a_read_cycle assignment, which is an e_assign
  assign mailbox_2_s1_in_a_read_cycle = (cpu_0_data_master_granted_mailbox_2_s1 & cpu_0_data_master_read) | (cpu_1_data_master_granted_mailbox_2_s1 & cpu_1_data_master_read) | (cpu_2_data_master_granted_mailbox_2_s1 & cpu_2_data_master_read) | (cpu_3_data_master_granted_mailbox_2_s1 & cpu_3_data_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = mailbox_2_s1_in_a_read_cycle;

  //mailbox_2_s1_waits_for_write in a cycle, which is an e_mux
  assign mailbox_2_s1_waits_for_write = mailbox_2_s1_in_a_write_cycle & 0;

  //mailbox_2_s1_in_a_write_cycle assignment, which is an e_assign
  assign mailbox_2_s1_in_a_write_cycle = (cpu_0_data_master_granted_mailbox_2_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_mailbox_2_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_mailbox_2_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_mailbox_2_s1 & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = mailbox_2_s1_in_a_write_cycle;

  assign wait_for_mailbox_2_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //mailbox_2/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_mailbox_2_s1 + cpu_1_data_master_granted_mailbox_2_s1 + cpu_2_data_master_granted_mailbox_2_s1 + cpu_3_data_master_granted_mailbox_2_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_mailbox_2_s1 + cpu_1_data_master_saved_grant_mailbox_2_s1 + cpu_2_data_master_saved_grant_mailbox_2_s1 + cpu_3_data_master_saved_grant_mailbox_2_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module mailbox_3_s1_arbitrator (
                                 // inputs:
                                  clk,
                                  cpu_0_data_master_address_to_slave,
                                  cpu_0_data_master_latency_counter,
                                  cpu_0_data_master_read,
                                  cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_0_data_master_write,
                                  cpu_0_data_master_writedata,
                                  cpu_1_data_master_address_to_slave,
                                  cpu_1_data_master_latency_counter,
                                  cpu_1_data_master_read,
                                  cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_1_data_master_write,
                                  cpu_1_data_master_writedata,
                                  cpu_2_data_master_address_to_slave,
                                  cpu_2_data_master_latency_counter,
                                  cpu_2_data_master_read,
                                  cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_2_data_master_write,
                                  cpu_2_data_master_writedata,
                                  cpu_3_data_master_address_to_slave,
                                  cpu_3_data_master_latency_counter,
                                  cpu_3_data_master_read,
                                  cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                  cpu_3_data_master_write,
                                  cpu_3_data_master_writedata,
                                  mailbox_3_s1_readdata,
                                  reset_n,

                                 // outputs:
                                  cpu_0_data_master_granted_mailbox_3_s1,
                                  cpu_0_data_master_qualified_request_mailbox_3_s1,
                                  cpu_0_data_master_read_data_valid_mailbox_3_s1,
                                  cpu_0_data_master_requests_mailbox_3_s1,
                                  cpu_1_data_master_granted_mailbox_3_s1,
                                  cpu_1_data_master_qualified_request_mailbox_3_s1,
                                  cpu_1_data_master_read_data_valid_mailbox_3_s1,
                                  cpu_1_data_master_requests_mailbox_3_s1,
                                  cpu_2_data_master_granted_mailbox_3_s1,
                                  cpu_2_data_master_qualified_request_mailbox_3_s1,
                                  cpu_2_data_master_read_data_valid_mailbox_3_s1,
                                  cpu_2_data_master_requests_mailbox_3_s1,
                                  cpu_3_data_master_granted_mailbox_3_s1,
                                  cpu_3_data_master_qualified_request_mailbox_3_s1,
                                  cpu_3_data_master_read_data_valid_mailbox_3_s1,
                                  cpu_3_data_master_requests_mailbox_3_s1,
                                  d1_mailbox_3_s1_end_xfer,
                                  mailbox_3_s1_address,
                                  mailbox_3_s1_chipselect,
                                  mailbox_3_s1_read,
                                  mailbox_3_s1_readdata_from_sa,
                                  mailbox_3_s1_reset_n,
                                  mailbox_3_s1_write,
                                  mailbox_3_s1_writedata
                               )
;

  output           cpu_0_data_master_granted_mailbox_3_s1;
  output           cpu_0_data_master_qualified_request_mailbox_3_s1;
  output           cpu_0_data_master_read_data_valid_mailbox_3_s1;
  output           cpu_0_data_master_requests_mailbox_3_s1;
  output           cpu_1_data_master_granted_mailbox_3_s1;
  output           cpu_1_data_master_qualified_request_mailbox_3_s1;
  output           cpu_1_data_master_read_data_valid_mailbox_3_s1;
  output           cpu_1_data_master_requests_mailbox_3_s1;
  output           cpu_2_data_master_granted_mailbox_3_s1;
  output           cpu_2_data_master_qualified_request_mailbox_3_s1;
  output           cpu_2_data_master_read_data_valid_mailbox_3_s1;
  output           cpu_2_data_master_requests_mailbox_3_s1;
  output           cpu_3_data_master_granted_mailbox_3_s1;
  output           cpu_3_data_master_qualified_request_mailbox_3_s1;
  output           cpu_3_data_master_read_data_valid_mailbox_3_s1;
  output           cpu_3_data_master_requests_mailbox_3_s1;
  output           d1_mailbox_3_s1_end_xfer;
  output  [  1: 0] mailbox_3_s1_address;
  output           mailbox_3_s1_chipselect;
  output           mailbox_3_s1_read;
  output  [ 31: 0] mailbox_3_s1_readdata_from_sa;
  output           mailbox_3_s1_reset_n;
  output           mailbox_3_s1_write;
  output  [ 31: 0] mailbox_3_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 31: 0] mailbox_3_s1_readdata;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_mailbox_3_s1;
  wire             cpu_0_data_master_qualified_request_mailbox_3_s1;
  wire             cpu_0_data_master_read_data_valid_mailbox_3_s1;
  wire             cpu_0_data_master_requests_mailbox_3_s1;
  wire             cpu_0_data_master_saved_grant_mailbox_3_s1;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_mailbox_3_s1;
  wire             cpu_1_data_master_qualified_request_mailbox_3_s1;
  wire             cpu_1_data_master_read_data_valid_mailbox_3_s1;
  wire             cpu_1_data_master_requests_mailbox_3_s1;
  wire             cpu_1_data_master_saved_grant_mailbox_3_s1;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_mailbox_3_s1;
  wire             cpu_2_data_master_qualified_request_mailbox_3_s1;
  wire             cpu_2_data_master_read_data_valid_mailbox_3_s1;
  wire             cpu_2_data_master_requests_mailbox_3_s1;
  wire             cpu_2_data_master_saved_grant_mailbox_3_s1;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_mailbox_3_s1;
  wire             cpu_3_data_master_qualified_request_mailbox_3_s1;
  wire             cpu_3_data_master_read_data_valid_mailbox_3_s1;
  wire             cpu_3_data_master_requests_mailbox_3_s1;
  wire             cpu_3_data_master_saved_grant_mailbox_3_s1;
  reg              d1_mailbox_3_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_mailbox_3_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_mailbox_3_s1;
  reg              last_cycle_cpu_1_data_master_granted_slave_mailbox_3_s1;
  reg              last_cycle_cpu_2_data_master_granted_slave_mailbox_3_s1;
  reg              last_cycle_cpu_3_data_master_granted_slave_mailbox_3_s1;
  wire    [  1: 0] mailbox_3_s1_address;
  wire             mailbox_3_s1_allgrants;
  wire             mailbox_3_s1_allow_new_arb_cycle;
  wire             mailbox_3_s1_any_bursting_master_saved_grant;
  wire             mailbox_3_s1_any_continuerequest;
  reg     [  3: 0] mailbox_3_s1_arb_addend;
  wire             mailbox_3_s1_arb_counter_enable;
  reg     [  2: 0] mailbox_3_s1_arb_share_counter;
  wire    [  2: 0] mailbox_3_s1_arb_share_counter_next_value;
  wire    [  2: 0] mailbox_3_s1_arb_share_set_values;
  wire    [  3: 0] mailbox_3_s1_arb_winner;
  wire             mailbox_3_s1_arbitration_holdoff_internal;
  wire             mailbox_3_s1_beginbursttransfer_internal;
  wire             mailbox_3_s1_begins_xfer;
  wire             mailbox_3_s1_chipselect;
  wire    [  7: 0] mailbox_3_s1_chosen_master_double_vector;
  wire    [  3: 0] mailbox_3_s1_chosen_master_rot_left;
  wire             mailbox_3_s1_end_xfer;
  wire             mailbox_3_s1_firsttransfer;
  wire    [  3: 0] mailbox_3_s1_grant_vector;
  wire             mailbox_3_s1_in_a_read_cycle;
  wire             mailbox_3_s1_in_a_write_cycle;
  wire    [  3: 0] mailbox_3_s1_master_qreq_vector;
  wire             mailbox_3_s1_non_bursting_master_requests;
  wire             mailbox_3_s1_read;
  wire    [ 31: 0] mailbox_3_s1_readdata_from_sa;
  reg              mailbox_3_s1_reg_firsttransfer;
  wire             mailbox_3_s1_reset_n;
  reg     [  3: 0] mailbox_3_s1_saved_chosen_master_vector;
  reg              mailbox_3_s1_slavearbiterlockenable;
  wire             mailbox_3_s1_slavearbiterlockenable2;
  wire             mailbox_3_s1_unreg_firsttransfer;
  wire             mailbox_3_s1_waits_for_read;
  wire             mailbox_3_s1_waits_for_write;
  wire             mailbox_3_s1_write;
  wire    [ 31: 0] mailbox_3_s1_writedata;
  wire    [ 24: 0] shifted_address_to_mailbox_3_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_3_s1_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_3_s1_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_mailbox_3_s1_from_cpu_3_data_master;
  wire             wait_for_mailbox_3_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~mailbox_3_s1_end_xfer;
    end


  assign mailbox_3_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_mailbox_3_s1 | cpu_1_data_master_qualified_request_mailbox_3_s1 | cpu_2_data_master_qualified_request_mailbox_3_s1 | cpu_3_data_master_qualified_request_mailbox_3_s1));
  //assign mailbox_3_s1_readdata_from_sa = mailbox_3_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign mailbox_3_s1_readdata_from_sa = mailbox_3_s1_readdata;

  assign cpu_0_data_master_requests_mailbox_3_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h80) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //mailbox_3_s1_arb_share_counter set values, which is an e_mux
  assign mailbox_3_s1_arb_share_set_values = 1;

  //mailbox_3_s1_non_bursting_master_requests mux, which is an e_mux
  assign mailbox_3_s1_non_bursting_master_requests = cpu_0_data_master_requests_mailbox_3_s1 |
    cpu_1_data_master_requests_mailbox_3_s1 |
    cpu_2_data_master_requests_mailbox_3_s1 |
    cpu_3_data_master_requests_mailbox_3_s1 |
    cpu_0_data_master_requests_mailbox_3_s1 |
    cpu_1_data_master_requests_mailbox_3_s1 |
    cpu_2_data_master_requests_mailbox_3_s1 |
    cpu_3_data_master_requests_mailbox_3_s1 |
    cpu_0_data_master_requests_mailbox_3_s1 |
    cpu_1_data_master_requests_mailbox_3_s1 |
    cpu_2_data_master_requests_mailbox_3_s1 |
    cpu_3_data_master_requests_mailbox_3_s1 |
    cpu_0_data_master_requests_mailbox_3_s1 |
    cpu_1_data_master_requests_mailbox_3_s1 |
    cpu_2_data_master_requests_mailbox_3_s1 |
    cpu_3_data_master_requests_mailbox_3_s1;

  //mailbox_3_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign mailbox_3_s1_any_bursting_master_saved_grant = 0;

  //mailbox_3_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign mailbox_3_s1_arb_share_counter_next_value = mailbox_3_s1_firsttransfer ? (mailbox_3_s1_arb_share_set_values - 1) : |mailbox_3_s1_arb_share_counter ? (mailbox_3_s1_arb_share_counter - 1) : 0;

  //mailbox_3_s1_allgrants all slave grants, which is an e_mux
  assign mailbox_3_s1_allgrants = (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector) |
    (|mailbox_3_s1_grant_vector);

  //mailbox_3_s1_end_xfer assignment, which is an e_assign
  assign mailbox_3_s1_end_xfer = ~(mailbox_3_s1_waits_for_read | mailbox_3_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_mailbox_3_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_mailbox_3_s1 = mailbox_3_s1_end_xfer & (~mailbox_3_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //mailbox_3_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign mailbox_3_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_mailbox_3_s1 & mailbox_3_s1_allgrants) | (end_xfer_arb_share_counter_term_mailbox_3_s1 & ~mailbox_3_s1_non_bursting_master_requests);

  //mailbox_3_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_3_s1_arb_share_counter <= 0;
      else if (mailbox_3_s1_arb_counter_enable)
          mailbox_3_s1_arb_share_counter <= mailbox_3_s1_arb_share_counter_next_value;
    end


  //mailbox_3_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_3_s1_slavearbiterlockenable <= 0;
      else if ((|mailbox_3_s1_master_qreq_vector & end_xfer_arb_share_counter_term_mailbox_3_s1) | (end_xfer_arb_share_counter_term_mailbox_3_s1 & ~mailbox_3_s1_non_bursting_master_requests))
          mailbox_3_s1_slavearbiterlockenable <= |mailbox_3_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master mailbox_3/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = mailbox_3_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //mailbox_3_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign mailbox_3_s1_slavearbiterlockenable2 = |mailbox_3_s1_arb_share_counter_next_value;

  //cpu_0/data_master mailbox_3/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = mailbox_3_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_1/data_master mailbox_3/s1 arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = mailbox_3_s1_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master mailbox_3/s1 arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = mailbox_3_s1_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted mailbox_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_mailbox_3_s1 <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_mailbox_3_s1 <= cpu_1_data_master_saved_grant_mailbox_3_s1 ? 1 : (mailbox_3_s1_arbitration_holdoff_internal | ~cpu_1_data_master_requests_mailbox_3_s1) ? 0 : last_cycle_cpu_1_data_master_granted_slave_mailbox_3_s1;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_mailbox_3_s1 & cpu_1_data_master_requests_mailbox_3_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_mailbox_3_s1 & cpu_1_data_master_requests_mailbox_3_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_mailbox_3_s1 & cpu_1_data_master_requests_mailbox_3_s1);

  //mailbox_3_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign mailbox_3_s1_any_continuerequest = cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest;

  //cpu_2/data_master mailbox_3/s1 arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = mailbox_3_s1_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master mailbox_3/s1 arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = mailbox_3_s1_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted mailbox_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_mailbox_3_s1 <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_mailbox_3_s1 <= cpu_2_data_master_saved_grant_mailbox_3_s1 ? 1 : (mailbox_3_s1_arbitration_holdoff_internal | ~cpu_2_data_master_requests_mailbox_3_s1) ? 0 : last_cycle_cpu_2_data_master_granted_slave_mailbox_3_s1;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_mailbox_3_s1 & cpu_2_data_master_requests_mailbox_3_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_mailbox_3_s1 & cpu_2_data_master_requests_mailbox_3_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_mailbox_3_s1 & cpu_2_data_master_requests_mailbox_3_s1);

  //cpu_3/data_master mailbox_3/s1 arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = mailbox_3_s1_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master mailbox_3/s1 arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = mailbox_3_s1_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted mailbox_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_mailbox_3_s1 <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_mailbox_3_s1 <= cpu_3_data_master_saved_grant_mailbox_3_s1 ? 1 : (mailbox_3_s1_arbitration_holdoff_internal | ~cpu_3_data_master_requests_mailbox_3_s1) ? 0 : last_cycle_cpu_3_data_master_granted_slave_mailbox_3_s1;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_mailbox_3_s1 & cpu_3_data_master_requests_mailbox_3_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_mailbox_3_s1 & cpu_3_data_master_requests_mailbox_3_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_mailbox_3_s1 & cpu_3_data_master_requests_mailbox_3_s1);

  assign cpu_0_data_master_qualified_request_mailbox_3_s1 = cpu_0_data_master_requests_mailbox_3_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_mailbox_3_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_mailbox_3_s1 = cpu_0_data_master_granted_mailbox_3_s1 & cpu_0_data_master_read & ~mailbox_3_s1_waits_for_read;

  //mailbox_3_s1_writedata mux, which is an e_mux
  assign mailbox_3_s1_writedata = (cpu_0_data_master_granted_mailbox_3_s1)? cpu_0_data_master_writedata :
    (cpu_1_data_master_granted_mailbox_3_s1)? cpu_1_data_master_writedata :
    (cpu_2_data_master_granted_mailbox_3_s1)? cpu_2_data_master_writedata :
    cpu_3_data_master_writedata;

  assign cpu_1_data_master_requests_mailbox_3_s1 = ({cpu_1_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h80) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //cpu_0/data_master granted mailbox_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_mailbox_3_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_mailbox_3_s1 <= cpu_0_data_master_saved_grant_mailbox_3_s1 ? 1 : (mailbox_3_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_mailbox_3_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_mailbox_3_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_mailbox_3_s1 & cpu_0_data_master_requests_mailbox_3_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_mailbox_3_s1 & cpu_0_data_master_requests_mailbox_3_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_mailbox_3_s1 & cpu_0_data_master_requests_mailbox_3_s1);

  assign cpu_1_data_master_qualified_request_mailbox_3_s1 = cpu_1_data_master_requests_mailbox_3_s1 & ~((cpu_1_data_master_read & ((cpu_1_data_master_latency_counter != 0) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_1_data_master_read_data_valid_mailbox_3_s1, which is an e_mux
  assign cpu_1_data_master_read_data_valid_mailbox_3_s1 = cpu_1_data_master_granted_mailbox_3_s1 & cpu_1_data_master_read & ~mailbox_3_s1_waits_for_read;

  assign cpu_2_data_master_requests_mailbox_3_s1 = ({cpu_2_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h80) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_mailbox_3_s1 = cpu_2_data_master_requests_mailbox_3_s1 & ~((cpu_2_data_master_read & ((cpu_2_data_master_latency_counter != 0) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_2_data_master_read_data_valid_mailbox_3_s1, which is an e_mux
  assign cpu_2_data_master_read_data_valid_mailbox_3_s1 = cpu_2_data_master_granted_mailbox_3_s1 & cpu_2_data_master_read & ~mailbox_3_s1_waits_for_read;

  assign cpu_3_data_master_requests_mailbox_3_s1 = ({cpu_3_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h80) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_mailbox_3_s1 = cpu_3_data_master_requests_mailbox_3_s1 & ~((cpu_3_data_master_read & ((cpu_3_data_master_latency_counter != 0) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock);
  //local readdatavalid cpu_3_data_master_read_data_valid_mailbox_3_s1, which is an e_mux
  assign cpu_3_data_master_read_data_valid_mailbox_3_s1 = cpu_3_data_master_granted_mailbox_3_s1 & cpu_3_data_master_read & ~mailbox_3_s1_waits_for_read;

  //allow new arb cycle for mailbox_3/s1, which is an e_assign
  assign mailbox_3_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_3_data_master_arbiterlock;

  //cpu_3/data_master assignment into master qualified-requests vector for mailbox_3/s1, which is an e_assign
  assign mailbox_3_s1_master_qreq_vector[0] = cpu_3_data_master_qualified_request_mailbox_3_s1;

  //cpu_3/data_master grant mailbox_3/s1, which is an e_assign
  assign cpu_3_data_master_granted_mailbox_3_s1 = mailbox_3_s1_grant_vector[0];

  //cpu_3/data_master saved-grant mailbox_3/s1, which is an e_assign
  assign cpu_3_data_master_saved_grant_mailbox_3_s1 = mailbox_3_s1_arb_winner[0] && cpu_3_data_master_requests_mailbox_3_s1;

  //cpu_2/data_master assignment into master qualified-requests vector for mailbox_3/s1, which is an e_assign
  assign mailbox_3_s1_master_qreq_vector[1] = cpu_2_data_master_qualified_request_mailbox_3_s1;

  //cpu_2/data_master grant mailbox_3/s1, which is an e_assign
  assign cpu_2_data_master_granted_mailbox_3_s1 = mailbox_3_s1_grant_vector[1];

  //cpu_2/data_master saved-grant mailbox_3/s1, which is an e_assign
  assign cpu_2_data_master_saved_grant_mailbox_3_s1 = mailbox_3_s1_arb_winner[1] && cpu_2_data_master_requests_mailbox_3_s1;

  //cpu_1/data_master assignment into master qualified-requests vector for mailbox_3/s1, which is an e_assign
  assign mailbox_3_s1_master_qreq_vector[2] = cpu_1_data_master_qualified_request_mailbox_3_s1;

  //cpu_1/data_master grant mailbox_3/s1, which is an e_assign
  assign cpu_1_data_master_granted_mailbox_3_s1 = mailbox_3_s1_grant_vector[2];

  //cpu_1/data_master saved-grant mailbox_3/s1, which is an e_assign
  assign cpu_1_data_master_saved_grant_mailbox_3_s1 = mailbox_3_s1_arb_winner[2] && cpu_1_data_master_requests_mailbox_3_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for mailbox_3/s1, which is an e_assign
  assign mailbox_3_s1_master_qreq_vector[3] = cpu_0_data_master_qualified_request_mailbox_3_s1;

  //cpu_0/data_master grant mailbox_3/s1, which is an e_assign
  assign cpu_0_data_master_granted_mailbox_3_s1 = mailbox_3_s1_grant_vector[3];

  //cpu_0/data_master saved-grant mailbox_3/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_mailbox_3_s1 = mailbox_3_s1_arb_winner[3] && cpu_0_data_master_requests_mailbox_3_s1;

  //mailbox_3/s1 chosen-master double-vector, which is an e_assign
  assign mailbox_3_s1_chosen_master_double_vector = {mailbox_3_s1_master_qreq_vector, mailbox_3_s1_master_qreq_vector} & ({~mailbox_3_s1_master_qreq_vector, ~mailbox_3_s1_master_qreq_vector} + mailbox_3_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign mailbox_3_s1_arb_winner = (mailbox_3_s1_allow_new_arb_cycle & | mailbox_3_s1_grant_vector) ? mailbox_3_s1_grant_vector : mailbox_3_s1_saved_chosen_master_vector;

  //saved mailbox_3_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_3_s1_saved_chosen_master_vector <= 0;
      else if (mailbox_3_s1_allow_new_arb_cycle)
          mailbox_3_s1_saved_chosen_master_vector <= |mailbox_3_s1_grant_vector ? mailbox_3_s1_grant_vector : mailbox_3_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign mailbox_3_s1_grant_vector = {(mailbox_3_s1_chosen_master_double_vector[3] | mailbox_3_s1_chosen_master_double_vector[7]),
    (mailbox_3_s1_chosen_master_double_vector[2] | mailbox_3_s1_chosen_master_double_vector[6]),
    (mailbox_3_s1_chosen_master_double_vector[1] | mailbox_3_s1_chosen_master_double_vector[5]),
    (mailbox_3_s1_chosen_master_double_vector[0] | mailbox_3_s1_chosen_master_double_vector[4])};

  //mailbox_3/s1 chosen master rotated left, which is an e_assign
  assign mailbox_3_s1_chosen_master_rot_left = (mailbox_3_s1_arb_winner << 1) ? (mailbox_3_s1_arb_winner << 1) : 1;

  //mailbox_3/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_3_s1_arb_addend <= 1;
      else if (|mailbox_3_s1_grant_vector)
          mailbox_3_s1_arb_addend <= mailbox_3_s1_end_xfer? mailbox_3_s1_chosen_master_rot_left : mailbox_3_s1_grant_vector;
    end


  //mailbox_3_s1_reset_n assignment, which is an e_assign
  assign mailbox_3_s1_reset_n = reset_n;

  assign mailbox_3_s1_chipselect = cpu_0_data_master_granted_mailbox_3_s1 | cpu_1_data_master_granted_mailbox_3_s1 | cpu_2_data_master_granted_mailbox_3_s1 | cpu_3_data_master_granted_mailbox_3_s1;
  //mailbox_3_s1_firsttransfer first transaction, which is an e_assign
  assign mailbox_3_s1_firsttransfer = mailbox_3_s1_begins_xfer ? mailbox_3_s1_unreg_firsttransfer : mailbox_3_s1_reg_firsttransfer;

  //mailbox_3_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign mailbox_3_s1_unreg_firsttransfer = ~(mailbox_3_s1_slavearbiterlockenable & mailbox_3_s1_any_continuerequest);

  //mailbox_3_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          mailbox_3_s1_reg_firsttransfer <= 1'b1;
      else if (mailbox_3_s1_begins_xfer)
          mailbox_3_s1_reg_firsttransfer <= mailbox_3_s1_unreg_firsttransfer;
    end


  //mailbox_3_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign mailbox_3_s1_beginbursttransfer_internal = mailbox_3_s1_begins_xfer;

  //mailbox_3_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign mailbox_3_s1_arbitration_holdoff_internal = mailbox_3_s1_begins_xfer & mailbox_3_s1_firsttransfer;

  //mailbox_3_s1_read assignment, which is an e_mux
  assign mailbox_3_s1_read = (cpu_0_data_master_granted_mailbox_3_s1 & cpu_0_data_master_read) | (cpu_1_data_master_granted_mailbox_3_s1 & cpu_1_data_master_read) | (cpu_2_data_master_granted_mailbox_3_s1 & cpu_2_data_master_read) | (cpu_3_data_master_granted_mailbox_3_s1 & cpu_3_data_master_read);

  //mailbox_3_s1_write assignment, which is an e_mux
  assign mailbox_3_s1_write = (cpu_0_data_master_granted_mailbox_3_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_mailbox_3_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_mailbox_3_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_mailbox_3_s1 & cpu_3_data_master_write);

  assign shifted_address_to_mailbox_3_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //mailbox_3_s1_address mux, which is an e_mux
  assign mailbox_3_s1_address = (cpu_0_data_master_granted_mailbox_3_s1)? (shifted_address_to_mailbox_3_s1_from_cpu_0_data_master >> 2) :
    (cpu_1_data_master_granted_mailbox_3_s1)? (shifted_address_to_mailbox_3_s1_from_cpu_1_data_master >> 2) :
    (cpu_2_data_master_granted_mailbox_3_s1)? (shifted_address_to_mailbox_3_s1_from_cpu_2_data_master >> 2) :
    (shifted_address_to_mailbox_3_s1_from_cpu_3_data_master >> 2);

  assign shifted_address_to_mailbox_3_s1_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_mailbox_3_s1_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_mailbox_3_s1_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  //d1_mailbox_3_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_mailbox_3_s1_end_xfer <= 1;
      else 
        d1_mailbox_3_s1_end_xfer <= mailbox_3_s1_end_xfer;
    end


  //mailbox_3_s1_waits_for_read in a cycle, which is an e_mux
  assign mailbox_3_s1_waits_for_read = mailbox_3_s1_in_a_read_cycle & mailbox_3_s1_begins_xfer;

  //mailbox_3_s1_in_a_read_cycle assignment, which is an e_assign
  assign mailbox_3_s1_in_a_read_cycle = (cpu_0_data_master_granted_mailbox_3_s1 & cpu_0_data_master_read) | (cpu_1_data_master_granted_mailbox_3_s1 & cpu_1_data_master_read) | (cpu_2_data_master_granted_mailbox_3_s1 & cpu_2_data_master_read) | (cpu_3_data_master_granted_mailbox_3_s1 & cpu_3_data_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = mailbox_3_s1_in_a_read_cycle;

  //mailbox_3_s1_waits_for_write in a cycle, which is an e_mux
  assign mailbox_3_s1_waits_for_write = mailbox_3_s1_in_a_write_cycle & 0;

  //mailbox_3_s1_in_a_write_cycle assignment, which is an e_assign
  assign mailbox_3_s1_in_a_write_cycle = (cpu_0_data_master_granted_mailbox_3_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_mailbox_3_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_mailbox_3_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_mailbox_3_s1 & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = mailbox_3_s1_in_a_write_cycle;

  assign wait_for_mailbox_3_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //mailbox_3/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_mailbox_3_s1 + cpu_1_data_master_granted_mailbox_3_s1 + cpu_2_data_master_granted_mailbox_3_s1 + cpu_3_data_master_granted_mailbox_3_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_mailbox_3_s1 + cpu_1_data_master_saved_grant_mailbox_3_s1 + cpu_2_data_master_saved_grant_mailbox_3_s1 + cpu_3_data_master_saved_grant_mailbox_3_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_0_in_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_1_instruction_master_address_to_slave,
                                            cpu_1_instruction_master_dbs_address,
                                            cpu_1_instruction_master_latency_counter,
                                            cpu_1_instruction_master_read,
                                            cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                            nios_system_clock_0_in_endofpacket,
                                            nios_system_clock_0_in_readdata,
                                            nios_system_clock_0_in_waitrequest,
                                            reset_n,

                                           // outputs:
                                            cpu_1_instruction_master_granted_nios_system_clock_0_in,
                                            cpu_1_instruction_master_qualified_request_nios_system_clock_0_in,
                                            cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in,
                                            cpu_1_instruction_master_requests_nios_system_clock_0_in,
                                            d1_nios_system_clock_0_in_end_xfer,
                                            nios_system_clock_0_in_address,
                                            nios_system_clock_0_in_byteenable,
                                            nios_system_clock_0_in_endofpacket_from_sa,
                                            nios_system_clock_0_in_nativeaddress,
                                            nios_system_clock_0_in_read,
                                            nios_system_clock_0_in_readdata_from_sa,
                                            nios_system_clock_0_in_reset_n,
                                            nios_system_clock_0_in_waitrequest_from_sa,
                                            nios_system_clock_0_in_write
                                         )
;

  output           cpu_1_instruction_master_granted_nios_system_clock_0_in;
  output           cpu_1_instruction_master_qualified_request_nios_system_clock_0_in;
  output           cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in;
  output           cpu_1_instruction_master_requests_nios_system_clock_0_in;
  output           d1_nios_system_clock_0_in_end_xfer;
  output  [ 22: 0] nios_system_clock_0_in_address;
  output  [  1: 0] nios_system_clock_0_in_byteenable;
  output           nios_system_clock_0_in_endofpacket_from_sa;
  output  [ 21: 0] nios_system_clock_0_in_nativeaddress;
  output           nios_system_clock_0_in_read;
  output  [ 15: 0] nios_system_clock_0_in_readdata_from_sa;
  output           nios_system_clock_0_in_reset_n;
  output           nios_system_clock_0_in_waitrequest_from_sa;
  output           nios_system_clock_0_in_write;
  input            clk;
  input   [ 24: 0] cpu_1_instruction_master_address_to_slave;
  input   [  1: 0] cpu_1_instruction_master_dbs_address;
  input            cpu_1_instruction_master_latency_counter;
  input            cpu_1_instruction_master_read;
  input            cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            nios_system_clock_0_in_endofpacket;
  input   [ 15: 0] nios_system_clock_0_in_readdata;
  input            nios_system_clock_0_in_waitrequest;
  input            reset_n;

  wire             cpu_1_instruction_master_arbiterlock;
  wire             cpu_1_instruction_master_arbiterlock2;
  wire             cpu_1_instruction_master_continuerequest;
  wire             cpu_1_instruction_master_granted_nios_system_clock_0_in;
  wire             cpu_1_instruction_master_qualified_request_nios_system_clock_0_in;
  wire             cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in;
  wire             cpu_1_instruction_master_requests_nios_system_clock_0_in;
  wire             cpu_1_instruction_master_saved_grant_nios_system_clock_0_in;
  reg              d1_nios_system_clock_0_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_0_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 22: 0] nios_system_clock_0_in_address;
  wire             nios_system_clock_0_in_allgrants;
  wire             nios_system_clock_0_in_allow_new_arb_cycle;
  wire             nios_system_clock_0_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_0_in_any_continuerequest;
  wire             nios_system_clock_0_in_arb_counter_enable;
  reg     [  1: 0] nios_system_clock_0_in_arb_share_counter;
  wire    [  1: 0] nios_system_clock_0_in_arb_share_counter_next_value;
  wire    [  1: 0] nios_system_clock_0_in_arb_share_set_values;
  wire             nios_system_clock_0_in_beginbursttransfer_internal;
  wire             nios_system_clock_0_in_begins_xfer;
  wire    [  1: 0] nios_system_clock_0_in_byteenable;
  wire             nios_system_clock_0_in_end_xfer;
  wire             nios_system_clock_0_in_endofpacket_from_sa;
  wire             nios_system_clock_0_in_firsttransfer;
  wire             nios_system_clock_0_in_grant_vector;
  wire             nios_system_clock_0_in_in_a_read_cycle;
  wire             nios_system_clock_0_in_in_a_write_cycle;
  wire             nios_system_clock_0_in_master_qreq_vector;
  wire    [ 21: 0] nios_system_clock_0_in_nativeaddress;
  wire             nios_system_clock_0_in_non_bursting_master_requests;
  wire             nios_system_clock_0_in_read;
  wire    [ 15: 0] nios_system_clock_0_in_readdata_from_sa;
  reg              nios_system_clock_0_in_reg_firsttransfer;
  wire             nios_system_clock_0_in_reset_n;
  reg              nios_system_clock_0_in_slavearbiterlockenable;
  wire             nios_system_clock_0_in_slavearbiterlockenable2;
  wire             nios_system_clock_0_in_unreg_firsttransfer;
  wire             nios_system_clock_0_in_waitrequest_from_sa;
  wire             nios_system_clock_0_in_waits_for_read;
  wire             nios_system_clock_0_in_waits_for_write;
  wire             nios_system_clock_0_in_write;
  wire             wait_for_nios_system_clock_0_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_0_in_end_xfer;
    end


  assign nios_system_clock_0_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_1_instruction_master_qualified_request_nios_system_clock_0_in));
  //assign nios_system_clock_0_in_readdata_from_sa = nios_system_clock_0_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_0_in_readdata_from_sa = nios_system_clock_0_in_readdata;

  assign cpu_1_instruction_master_requests_nios_system_clock_0_in = (({cpu_1_instruction_master_address_to_slave[24 : 23] , 23'b0} == 25'h800000) & (cpu_1_instruction_master_read)) & cpu_1_instruction_master_read;
  //assign nios_system_clock_0_in_waitrequest_from_sa = nios_system_clock_0_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_0_in_waitrequest_from_sa = nios_system_clock_0_in_waitrequest;

  //nios_system_clock_0_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_0_in_arb_share_set_values = (cpu_1_instruction_master_granted_nios_system_clock_0_in)? 2 :
    1;

  //nios_system_clock_0_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_0_in_non_bursting_master_requests = cpu_1_instruction_master_requests_nios_system_clock_0_in;

  //nios_system_clock_0_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_0_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_0_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_0_in_arb_share_counter_next_value = nios_system_clock_0_in_firsttransfer ? (nios_system_clock_0_in_arb_share_set_values - 1) : |nios_system_clock_0_in_arb_share_counter ? (nios_system_clock_0_in_arb_share_counter - 1) : 0;

  //nios_system_clock_0_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_0_in_allgrants = |nios_system_clock_0_in_grant_vector;

  //nios_system_clock_0_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_0_in_end_xfer = ~(nios_system_clock_0_in_waits_for_read | nios_system_clock_0_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_0_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_0_in = nios_system_clock_0_in_end_xfer & (~nios_system_clock_0_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_0_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_0_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_0_in & nios_system_clock_0_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_0_in & ~nios_system_clock_0_in_non_bursting_master_requests);

  //nios_system_clock_0_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_0_in_arb_share_counter <= 0;
      else if (nios_system_clock_0_in_arb_counter_enable)
          nios_system_clock_0_in_arb_share_counter <= nios_system_clock_0_in_arb_share_counter_next_value;
    end


  //nios_system_clock_0_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_0_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_0_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_0_in) | (end_xfer_arb_share_counter_term_nios_system_clock_0_in & ~nios_system_clock_0_in_non_bursting_master_requests))
          nios_system_clock_0_in_slavearbiterlockenable <= |nios_system_clock_0_in_arb_share_counter_next_value;
    end


  //cpu_1/instruction_master nios_system_clock_0/in arbiterlock, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock = nios_system_clock_0_in_slavearbiterlockenable & cpu_1_instruction_master_continuerequest;

  //nios_system_clock_0_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_0_in_slavearbiterlockenable2 = |nios_system_clock_0_in_arb_share_counter_next_value;

  //cpu_1/instruction_master nios_system_clock_0/in arbiterlock2, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock2 = nios_system_clock_0_in_slavearbiterlockenable2 & cpu_1_instruction_master_continuerequest;

  //nios_system_clock_0_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_0_in_any_continuerequest = 1;

  //cpu_1_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_1_instruction_master_continuerequest = 1;

  assign cpu_1_instruction_master_qualified_request_nios_system_clock_0_in = cpu_1_instruction_master_requests_nios_system_clock_0_in & ~((cpu_1_instruction_master_read & ((cpu_1_instruction_master_latency_counter != 0) | (|cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))));
  //local readdatavalid cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in, which is an e_mux
  assign cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in = cpu_1_instruction_master_granted_nios_system_clock_0_in & cpu_1_instruction_master_read & ~nios_system_clock_0_in_waits_for_read;

  //assign nios_system_clock_0_in_endofpacket_from_sa = nios_system_clock_0_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_0_in_endofpacket_from_sa = nios_system_clock_0_in_endofpacket;

  //master is always granted when requested
  assign cpu_1_instruction_master_granted_nios_system_clock_0_in = cpu_1_instruction_master_qualified_request_nios_system_clock_0_in;

  //cpu_1/instruction_master saved-grant nios_system_clock_0/in, which is an e_assign
  assign cpu_1_instruction_master_saved_grant_nios_system_clock_0_in = cpu_1_instruction_master_requests_nios_system_clock_0_in;

  //allow new arb cycle for nios_system_clock_0/in, which is an e_assign
  assign nios_system_clock_0_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_0_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_0_in_master_qreq_vector = 1;

  //nios_system_clock_0_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_0_in_reset_n = reset_n;

  //nios_system_clock_0_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_0_in_firsttransfer = nios_system_clock_0_in_begins_xfer ? nios_system_clock_0_in_unreg_firsttransfer : nios_system_clock_0_in_reg_firsttransfer;

  //nios_system_clock_0_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_0_in_unreg_firsttransfer = ~(nios_system_clock_0_in_slavearbiterlockenable & nios_system_clock_0_in_any_continuerequest);

  //nios_system_clock_0_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_0_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_0_in_begins_xfer)
          nios_system_clock_0_in_reg_firsttransfer <= nios_system_clock_0_in_unreg_firsttransfer;
    end


  //nios_system_clock_0_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_0_in_beginbursttransfer_internal = nios_system_clock_0_in_begins_xfer;

  //nios_system_clock_0_in_read assignment, which is an e_mux
  assign nios_system_clock_0_in_read = cpu_1_instruction_master_granted_nios_system_clock_0_in & cpu_1_instruction_master_read;

  //nios_system_clock_0_in_write assignment, which is an e_mux
  assign nios_system_clock_0_in_write = 0;

  //nios_system_clock_0_in_address mux, which is an e_mux
  assign nios_system_clock_0_in_address = {cpu_1_instruction_master_address_to_slave >> 2,
    cpu_1_instruction_master_dbs_address[1],
    {1 {1'b0}}};

  //slaveid nios_system_clock_0_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_0_in_nativeaddress = cpu_1_instruction_master_address_to_slave >> 2;

  //d1_nios_system_clock_0_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_0_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_0_in_end_xfer <= nios_system_clock_0_in_end_xfer;
    end


  //nios_system_clock_0_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_0_in_waits_for_read = nios_system_clock_0_in_in_a_read_cycle & nios_system_clock_0_in_waitrequest_from_sa;

  //nios_system_clock_0_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_0_in_in_a_read_cycle = cpu_1_instruction_master_granted_nios_system_clock_0_in & cpu_1_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_0_in_in_a_read_cycle;

  //nios_system_clock_0_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_0_in_waits_for_write = nios_system_clock_0_in_in_a_write_cycle & nios_system_clock_0_in_waitrequest_from_sa;

  //nios_system_clock_0_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_0_in_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_0_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_0_in_counter = 0;
  //nios_system_clock_0_in_byteenable byte enable port mux, which is an e_mux
  assign nios_system_clock_0_in_byteenable = -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_0/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_0_out_arbitrator (
                                            // inputs:
                                             clk,
                                             d1_sdram_0_s1_end_xfer,
                                             nios_system_clock_0_out_address,
                                             nios_system_clock_0_out_byteenable,
                                             nios_system_clock_0_out_granted_sdram_0_s1,
                                             nios_system_clock_0_out_qualified_request_sdram_0_s1,
                                             nios_system_clock_0_out_read,
                                             nios_system_clock_0_out_read_data_valid_sdram_0_s1,
                                             nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register,
                                             nios_system_clock_0_out_requests_sdram_0_s1,
                                             nios_system_clock_0_out_write,
                                             nios_system_clock_0_out_writedata,
                                             reset_n,
                                             sdram_0_s1_readdata_from_sa,
                                             sdram_0_s1_waitrequest_from_sa,

                                            // outputs:
                                             nios_system_clock_0_out_address_to_slave,
                                             nios_system_clock_0_out_readdata,
                                             nios_system_clock_0_out_reset_n,
                                             nios_system_clock_0_out_waitrequest
                                          )
;

  output  [ 22: 0] nios_system_clock_0_out_address_to_slave;
  output  [ 15: 0] nios_system_clock_0_out_readdata;
  output           nios_system_clock_0_out_reset_n;
  output           nios_system_clock_0_out_waitrequest;
  input            clk;
  input            d1_sdram_0_s1_end_xfer;
  input   [ 22: 0] nios_system_clock_0_out_address;
  input   [  1: 0] nios_system_clock_0_out_byteenable;
  input            nios_system_clock_0_out_granted_sdram_0_s1;
  input            nios_system_clock_0_out_qualified_request_sdram_0_s1;
  input            nios_system_clock_0_out_read;
  input            nios_system_clock_0_out_read_data_valid_sdram_0_s1;
  input            nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register;
  input            nios_system_clock_0_out_requests_sdram_0_s1;
  input            nios_system_clock_0_out_write;
  input   [ 15: 0] nios_system_clock_0_out_writedata;
  input            reset_n;
  input   [ 15: 0] sdram_0_s1_readdata_from_sa;
  input            sdram_0_s1_waitrequest_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 22: 0] nios_system_clock_0_out_address_last_time;
  wire    [ 22: 0] nios_system_clock_0_out_address_to_slave;
  reg     [  1: 0] nios_system_clock_0_out_byteenable_last_time;
  reg              nios_system_clock_0_out_read_last_time;
  wire    [ 15: 0] nios_system_clock_0_out_readdata;
  wire             nios_system_clock_0_out_reset_n;
  wire             nios_system_clock_0_out_run;
  wire             nios_system_clock_0_out_waitrequest;
  reg              nios_system_clock_0_out_write_last_time;
  reg     [ 15: 0] nios_system_clock_0_out_writedata_last_time;
  wire             r_3;
  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (nios_system_clock_0_out_qualified_request_sdram_0_s1 | nios_system_clock_0_out_read_data_valid_sdram_0_s1 | ~nios_system_clock_0_out_requests_sdram_0_s1) & (nios_system_clock_0_out_granted_sdram_0_s1 | ~nios_system_clock_0_out_qualified_request_sdram_0_s1) & ((~nios_system_clock_0_out_qualified_request_sdram_0_s1 | ~nios_system_clock_0_out_read | (nios_system_clock_0_out_read_data_valid_sdram_0_s1 & nios_system_clock_0_out_read))) & ((~nios_system_clock_0_out_qualified_request_sdram_0_s1 | ~(nios_system_clock_0_out_read | nios_system_clock_0_out_write) | (1 & ~sdram_0_s1_waitrequest_from_sa & (nios_system_clock_0_out_read | nios_system_clock_0_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_0_out_run = r_3;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_0_out_address_to_slave = nios_system_clock_0_out_address;

  //nios_system_clock_0/out readdata mux, which is an e_mux
  assign nios_system_clock_0_out_readdata = sdram_0_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_0_out_waitrequest = ~nios_system_clock_0_out_run;

  //nios_system_clock_0_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_0_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_0_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_0_out_address_last_time <= 0;
      else 
        nios_system_clock_0_out_address_last_time <= nios_system_clock_0_out_address;
    end


  //nios_system_clock_0/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_0_out_waitrequest & (nios_system_clock_0_out_read | nios_system_clock_0_out_write);
    end


  //nios_system_clock_0_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_0_out_address != nios_system_clock_0_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_0_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_0_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_0_out_byteenable_last_time <= 0;
      else 
        nios_system_clock_0_out_byteenable_last_time <= nios_system_clock_0_out_byteenable;
    end


  //nios_system_clock_0_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_0_out_byteenable != nios_system_clock_0_out_byteenable_last_time))
        begin
          $write("%0d ns: nios_system_clock_0_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_0_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_0_out_read_last_time <= 0;
      else 
        nios_system_clock_0_out_read_last_time <= nios_system_clock_0_out_read;
    end


  //nios_system_clock_0_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_0_out_read != nios_system_clock_0_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_0_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_0_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_0_out_write_last_time <= 0;
      else 
        nios_system_clock_0_out_write_last_time <= nios_system_clock_0_out_write;
    end


  //nios_system_clock_0_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_0_out_write != nios_system_clock_0_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_0_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_0_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_0_out_writedata_last_time <= 0;
      else 
        nios_system_clock_0_out_writedata_last_time <= nios_system_clock_0_out_writedata;
    end


  //nios_system_clock_0_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_0_out_writedata != nios_system_clock_0_out_writedata_last_time) & nios_system_clock_0_out_write)
        begin
          $write("%0d ns: nios_system_clock_0_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_1_in_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_1_data_master_address_to_slave,
                                            cpu_1_data_master_byteenable,
                                            cpu_1_data_master_dbs_address,
                                            cpu_1_data_master_dbs_write_16,
                                            cpu_1_data_master_latency_counter,
                                            cpu_1_data_master_read,
                                            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                            cpu_1_data_master_write,
                                            nios_system_clock_1_in_endofpacket,
                                            nios_system_clock_1_in_readdata,
                                            nios_system_clock_1_in_waitrequest,
                                            reset_n,

                                           // outputs:
                                            cpu_1_data_master_byteenable_nios_system_clock_1_in,
                                            cpu_1_data_master_granted_nios_system_clock_1_in,
                                            cpu_1_data_master_qualified_request_nios_system_clock_1_in,
                                            cpu_1_data_master_read_data_valid_nios_system_clock_1_in,
                                            cpu_1_data_master_requests_nios_system_clock_1_in,
                                            d1_nios_system_clock_1_in_end_xfer,
                                            nios_system_clock_1_in_address,
                                            nios_system_clock_1_in_byteenable,
                                            nios_system_clock_1_in_endofpacket_from_sa,
                                            nios_system_clock_1_in_nativeaddress,
                                            nios_system_clock_1_in_read,
                                            nios_system_clock_1_in_readdata_from_sa,
                                            nios_system_clock_1_in_reset_n,
                                            nios_system_clock_1_in_waitrequest_from_sa,
                                            nios_system_clock_1_in_write,
                                            nios_system_clock_1_in_writedata
                                         )
;

  output  [  1: 0] cpu_1_data_master_byteenable_nios_system_clock_1_in;
  output           cpu_1_data_master_granted_nios_system_clock_1_in;
  output           cpu_1_data_master_qualified_request_nios_system_clock_1_in;
  output           cpu_1_data_master_read_data_valid_nios_system_clock_1_in;
  output           cpu_1_data_master_requests_nios_system_clock_1_in;
  output           d1_nios_system_clock_1_in_end_xfer;
  output  [ 22: 0] nios_system_clock_1_in_address;
  output  [  1: 0] nios_system_clock_1_in_byteenable;
  output           nios_system_clock_1_in_endofpacket_from_sa;
  output  [ 21: 0] nios_system_clock_1_in_nativeaddress;
  output           nios_system_clock_1_in_read;
  output  [ 15: 0] nios_system_clock_1_in_readdata_from_sa;
  output           nios_system_clock_1_in_reset_n;
  output           nios_system_clock_1_in_waitrequest_from_sa;
  output           nios_system_clock_1_in_write;
  output  [ 15: 0] nios_system_clock_1_in_writedata;
  input            clk;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input   [  3: 0] cpu_1_data_master_byteenable;
  input   [  1: 0] cpu_1_data_master_dbs_address;
  input   [ 15: 0] cpu_1_data_master_dbs_write_16;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input            nios_system_clock_1_in_endofpacket;
  input   [ 15: 0] nios_system_clock_1_in_readdata;
  input            nios_system_clock_1_in_waitrequest;
  input            reset_n;

  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire    [  1: 0] cpu_1_data_master_byteenable_nios_system_clock_1_in;
  wire    [  1: 0] cpu_1_data_master_byteenable_nios_system_clock_1_in_segment_0;
  wire    [  1: 0] cpu_1_data_master_byteenable_nios_system_clock_1_in_segment_1;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_nios_system_clock_1_in;
  wire             cpu_1_data_master_qualified_request_nios_system_clock_1_in;
  wire             cpu_1_data_master_read_data_valid_nios_system_clock_1_in;
  wire             cpu_1_data_master_requests_nios_system_clock_1_in;
  wire             cpu_1_data_master_saved_grant_nios_system_clock_1_in;
  reg              d1_nios_system_clock_1_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_1_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 22: 0] nios_system_clock_1_in_address;
  wire             nios_system_clock_1_in_allgrants;
  wire             nios_system_clock_1_in_allow_new_arb_cycle;
  wire             nios_system_clock_1_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_1_in_any_continuerequest;
  wire             nios_system_clock_1_in_arb_counter_enable;
  reg     [  2: 0] nios_system_clock_1_in_arb_share_counter;
  wire    [  2: 0] nios_system_clock_1_in_arb_share_counter_next_value;
  wire    [  2: 0] nios_system_clock_1_in_arb_share_set_values;
  wire             nios_system_clock_1_in_beginbursttransfer_internal;
  wire             nios_system_clock_1_in_begins_xfer;
  wire    [  1: 0] nios_system_clock_1_in_byteenable;
  wire             nios_system_clock_1_in_end_xfer;
  wire             nios_system_clock_1_in_endofpacket_from_sa;
  wire             nios_system_clock_1_in_firsttransfer;
  wire             nios_system_clock_1_in_grant_vector;
  wire             nios_system_clock_1_in_in_a_read_cycle;
  wire             nios_system_clock_1_in_in_a_write_cycle;
  wire             nios_system_clock_1_in_master_qreq_vector;
  wire    [ 21: 0] nios_system_clock_1_in_nativeaddress;
  wire             nios_system_clock_1_in_non_bursting_master_requests;
  wire             nios_system_clock_1_in_read;
  wire    [ 15: 0] nios_system_clock_1_in_readdata_from_sa;
  reg              nios_system_clock_1_in_reg_firsttransfer;
  wire             nios_system_clock_1_in_reset_n;
  reg              nios_system_clock_1_in_slavearbiterlockenable;
  wire             nios_system_clock_1_in_slavearbiterlockenable2;
  wire             nios_system_clock_1_in_unreg_firsttransfer;
  wire             nios_system_clock_1_in_waitrequest_from_sa;
  wire             nios_system_clock_1_in_waits_for_read;
  wire             nios_system_clock_1_in_waits_for_write;
  wire             nios_system_clock_1_in_write;
  wire    [ 15: 0] nios_system_clock_1_in_writedata;
  wire             wait_for_nios_system_clock_1_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_1_in_end_xfer;
    end


  assign nios_system_clock_1_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_1_data_master_qualified_request_nios_system_clock_1_in));
  //assign nios_system_clock_1_in_readdata_from_sa = nios_system_clock_1_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_1_in_readdata_from_sa = nios_system_clock_1_in_readdata;

  assign cpu_1_data_master_requests_nios_system_clock_1_in = ({cpu_1_data_master_address_to_slave[24 : 23] , 23'b0} == 25'h800000) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //assign nios_system_clock_1_in_waitrequest_from_sa = nios_system_clock_1_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_1_in_waitrequest_from_sa = nios_system_clock_1_in_waitrequest;

  //nios_system_clock_1_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_1_in_arb_share_set_values = (cpu_1_data_master_granted_nios_system_clock_1_in)? 2 :
    1;

  //nios_system_clock_1_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_1_in_non_bursting_master_requests = cpu_1_data_master_requests_nios_system_clock_1_in;

  //nios_system_clock_1_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_1_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_1_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_1_in_arb_share_counter_next_value = nios_system_clock_1_in_firsttransfer ? (nios_system_clock_1_in_arb_share_set_values - 1) : |nios_system_clock_1_in_arb_share_counter ? (nios_system_clock_1_in_arb_share_counter - 1) : 0;

  //nios_system_clock_1_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_1_in_allgrants = |nios_system_clock_1_in_grant_vector;

  //nios_system_clock_1_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_1_in_end_xfer = ~(nios_system_clock_1_in_waits_for_read | nios_system_clock_1_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_1_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_1_in = nios_system_clock_1_in_end_xfer & (~nios_system_clock_1_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_1_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_1_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_1_in & nios_system_clock_1_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_1_in & ~nios_system_clock_1_in_non_bursting_master_requests);

  //nios_system_clock_1_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_1_in_arb_share_counter <= 0;
      else if (nios_system_clock_1_in_arb_counter_enable)
          nios_system_clock_1_in_arb_share_counter <= nios_system_clock_1_in_arb_share_counter_next_value;
    end


  //nios_system_clock_1_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_1_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_1_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_1_in) | (end_xfer_arb_share_counter_term_nios_system_clock_1_in & ~nios_system_clock_1_in_non_bursting_master_requests))
          nios_system_clock_1_in_slavearbiterlockenable <= |nios_system_clock_1_in_arb_share_counter_next_value;
    end


  //cpu_1/data_master nios_system_clock_1/in arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = nios_system_clock_1_in_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //nios_system_clock_1_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_1_in_slavearbiterlockenable2 = |nios_system_clock_1_in_arb_share_counter_next_value;

  //cpu_1/data_master nios_system_clock_1/in arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = nios_system_clock_1_in_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //nios_system_clock_1_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_1_in_any_continuerequest = 1;

  //cpu_1_data_master_continuerequest continued request, which is an e_assign
  assign cpu_1_data_master_continuerequest = 1;

  assign cpu_1_data_master_qualified_request_nios_system_clock_1_in = cpu_1_data_master_requests_nios_system_clock_1_in & ~((cpu_1_data_master_read & ((cpu_1_data_master_latency_counter != 0) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | ((!cpu_1_data_master_byteenable_nios_system_clock_1_in) & cpu_1_data_master_write));
  //local readdatavalid cpu_1_data_master_read_data_valid_nios_system_clock_1_in, which is an e_mux
  assign cpu_1_data_master_read_data_valid_nios_system_clock_1_in = cpu_1_data_master_granted_nios_system_clock_1_in & cpu_1_data_master_read & ~nios_system_clock_1_in_waits_for_read;

  //nios_system_clock_1_in_writedata mux, which is an e_mux
  assign nios_system_clock_1_in_writedata = cpu_1_data_master_dbs_write_16;

  //assign nios_system_clock_1_in_endofpacket_from_sa = nios_system_clock_1_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_1_in_endofpacket_from_sa = nios_system_clock_1_in_endofpacket;

  //master is always granted when requested
  assign cpu_1_data_master_granted_nios_system_clock_1_in = cpu_1_data_master_qualified_request_nios_system_clock_1_in;

  //cpu_1/data_master saved-grant nios_system_clock_1/in, which is an e_assign
  assign cpu_1_data_master_saved_grant_nios_system_clock_1_in = cpu_1_data_master_requests_nios_system_clock_1_in;

  //allow new arb cycle for nios_system_clock_1/in, which is an e_assign
  assign nios_system_clock_1_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_1_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_1_in_master_qreq_vector = 1;

  //nios_system_clock_1_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_1_in_reset_n = reset_n;

  //nios_system_clock_1_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_1_in_firsttransfer = nios_system_clock_1_in_begins_xfer ? nios_system_clock_1_in_unreg_firsttransfer : nios_system_clock_1_in_reg_firsttransfer;

  //nios_system_clock_1_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_1_in_unreg_firsttransfer = ~(nios_system_clock_1_in_slavearbiterlockenable & nios_system_clock_1_in_any_continuerequest);

  //nios_system_clock_1_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_1_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_1_in_begins_xfer)
          nios_system_clock_1_in_reg_firsttransfer <= nios_system_clock_1_in_unreg_firsttransfer;
    end


  //nios_system_clock_1_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_1_in_beginbursttransfer_internal = nios_system_clock_1_in_begins_xfer;

  //nios_system_clock_1_in_read assignment, which is an e_mux
  assign nios_system_clock_1_in_read = cpu_1_data_master_granted_nios_system_clock_1_in & cpu_1_data_master_read;

  //nios_system_clock_1_in_write assignment, which is an e_mux
  assign nios_system_clock_1_in_write = cpu_1_data_master_granted_nios_system_clock_1_in & cpu_1_data_master_write;

  //nios_system_clock_1_in_address mux, which is an e_mux
  assign nios_system_clock_1_in_address = {cpu_1_data_master_address_to_slave >> 2,
    cpu_1_data_master_dbs_address[1],
    {1 {1'b0}}};

  //slaveid nios_system_clock_1_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_1_in_nativeaddress = cpu_1_data_master_address_to_slave >> 2;

  //d1_nios_system_clock_1_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_1_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_1_in_end_xfer <= nios_system_clock_1_in_end_xfer;
    end


  //nios_system_clock_1_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_1_in_waits_for_read = nios_system_clock_1_in_in_a_read_cycle & nios_system_clock_1_in_waitrequest_from_sa;

  //nios_system_clock_1_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_1_in_in_a_read_cycle = cpu_1_data_master_granted_nios_system_clock_1_in & cpu_1_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_1_in_in_a_read_cycle;

  //nios_system_clock_1_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_1_in_waits_for_write = nios_system_clock_1_in_in_a_write_cycle & nios_system_clock_1_in_waitrequest_from_sa;

  //nios_system_clock_1_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_1_in_in_a_write_cycle = cpu_1_data_master_granted_nios_system_clock_1_in & cpu_1_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_1_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_1_in_counter = 0;
  //nios_system_clock_1_in_byteenable byte enable port mux, which is an e_mux
  assign nios_system_clock_1_in_byteenable = (cpu_1_data_master_granted_nios_system_clock_1_in)? cpu_1_data_master_byteenable_nios_system_clock_1_in :
    -1;

  assign {cpu_1_data_master_byteenable_nios_system_clock_1_in_segment_1,
cpu_1_data_master_byteenable_nios_system_clock_1_in_segment_0} = cpu_1_data_master_byteenable;
  assign cpu_1_data_master_byteenable_nios_system_clock_1_in = ((cpu_1_data_master_dbs_address[1] == 0))? cpu_1_data_master_byteenable_nios_system_clock_1_in_segment_0 :
    cpu_1_data_master_byteenable_nios_system_clock_1_in_segment_1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_1/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_1_out_arbitrator (
                                            // inputs:
                                             clk,
                                             d1_sdram_0_s1_end_xfer,
                                             nios_system_clock_1_out_address,
                                             nios_system_clock_1_out_byteenable,
                                             nios_system_clock_1_out_granted_sdram_0_s1,
                                             nios_system_clock_1_out_qualified_request_sdram_0_s1,
                                             nios_system_clock_1_out_read,
                                             nios_system_clock_1_out_read_data_valid_sdram_0_s1,
                                             nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register,
                                             nios_system_clock_1_out_requests_sdram_0_s1,
                                             nios_system_clock_1_out_write,
                                             nios_system_clock_1_out_writedata,
                                             reset_n,
                                             sdram_0_s1_readdata_from_sa,
                                             sdram_0_s1_waitrequest_from_sa,

                                            // outputs:
                                             nios_system_clock_1_out_address_to_slave,
                                             nios_system_clock_1_out_readdata,
                                             nios_system_clock_1_out_reset_n,
                                             nios_system_clock_1_out_waitrequest
                                          )
;

  output  [ 22: 0] nios_system_clock_1_out_address_to_slave;
  output  [ 15: 0] nios_system_clock_1_out_readdata;
  output           nios_system_clock_1_out_reset_n;
  output           nios_system_clock_1_out_waitrequest;
  input            clk;
  input            d1_sdram_0_s1_end_xfer;
  input   [ 22: 0] nios_system_clock_1_out_address;
  input   [  1: 0] nios_system_clock_1_out_byteenable;
  input            nios_system_clock_1_out_granted_sdram_0_s1;
  input            nios_system_clock_1_out_qualified_request_sdram_0_s1;
  input            nios_system_clock_1_out_read;
  input            nios_system_clock_1_out_read_data_valid_sdram_0_s1;
  input            nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register;
  input            nios_system_clock_1_out_requests_sdram_0_s1;
  input            nios_system_clock_1_out_write;
  input   [ 15: 0] nios_system_clock_1_out_writedata;
  input            reset_n;
  input   [ 15: 0] sdram_0_s1_readdata_from_sa;
  input            sdram_0_s1_waitrequest_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 22: 0] nios_system_clock_1_out_address_last_time;
  wire    [ 22: 0] nios_system_clock_1_out_address_to_slave;
  reg     [  1: 0] nios_system_clock_1_out_byteenable_last_time;
  reg              nios_system_clock_1_out_read_last_time;
  wire    [ 15: 0] nios_system_clock_1_out_readdata;
  wire             nios_system_clock_1_out_reset_n;
  wire             nios_system_clock_1_out_run;
  wire             nios_system_clock_1_out_waitrequest;
  reg              nios_system_clock_1_out_write_last_time;
  reg     [ 15: 0] nios_system_clock_1_out_writedata_last_time;
  wire             r_3;
  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (nios_system_clock_1_out_qualified_request_sdram_0_s1 | nios_system_clock_1_out_read_data_valid_sdram_0_s1 | ~nios_system_clock_1_out_requests_sdram_0_s1) & (nios_system_clock_1_out_granted_sdram_0_s1 | ~nios_system_clock_1_out_qualified_request_sdram_0_s1) & ((~nios_system_clock_1_out_qualified_request_sdram_0_s1 | ~nios_system_clock_1_out_read | (nios_system_clock_1_out_read_data_valid_sdram_0_s1 & nios_system_clock_1_out_read))) & ((~nios_system_clock_1_out_qualified_request_sdram_0_s1 | ~(nios_system_clock_1_out_read | nios_system_clock_1_out_write) | (1 & ~sdram_0_s1_waitrequest_from_sa & (nios_system_clock_1_out_read | nios_system_clock_1_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_1_out_run = r_3;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_1_out_address_to_slave = nios_system_clock_1_out_address;

  //nios_system_clock_1/out readdata mux, which is an e_mux
  assign nios_system_clock_1_out_readdata = sdram_0_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_1_out_waitrequest = ~nios_system_clock_1_out_run;

  //nios_system_clock_1_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_1_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_1_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_1_out_address_last_time <= 0;
      else 
        nios_system_clock_1_out_address_last_time <= nios_system_clock_1_out_address;
    end


  //nios_system_clock_1/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_1_out_waitrequest & (nios_system_clock_1_out_read | nios_system_clock_1_out_write);
    end


  //nios_system_clock_1_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_1_out_address != nios_system_clock_1_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_1_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_1_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_1_out_byteenable_last_time <= 0;
      else 
        nios_system_clock_1_out_byteenable_last_time <= nios_system_clock_1_out_byteenable;
    end


  //nios_system_clock_1_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_1_out_byteenable != nios_system_clock_1_out_byteenable_last_time))
        begin
          $write("%0d ns: nios_system_clock_1_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_1_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_1_out_read_last_time <= 0;
      else 
        nios_system_clock_1_out_read_last_time <= nios_system_clock_1_out_read;
    end


  //nios_system_clock_1_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_1_out_read != nios_system_clock_1_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_1_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_1_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_1_out_write_last_time <= 0;
      else 
        nios_system_clock_1_out_write_last_time <= nios_system_clock_1_out_write;
    end


  //nios_system_clock_1_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_1_out_write != nios_system_clock_1_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_1_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_1_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_1_out_writedata_last_time <= 0;
      else 
        nios_system_clock_1_out_writedata_last_time <= nios_system_clock_1_out_writedata;
    end


  //nios_system_clock_1_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_1_out_writedata != nios_system_clock_1_out_writedata_last_time) & nios_system_clock_1_out_write)
        begin
          $write("%0d ns: nios_system_clock_1_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_10_in_arbitrator (
                                            // inputs:
                                             clk,
                                             cpu_2_data_master_address_to_slave,
                                             cpu_2_data_master_byteenable,
                                             cpu_2_data_master_dbs_address,
                                             cpu_2_data_master_dbs_write_8,
                                             cpu_2_data_master_latency_counter,
                                             cpu_2_data_master_read,
                                             cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                             cpu_2_data_master_write,
                                             nios_system_clock_10_in_endofpacket,
                                             nios_system_clock_10_in_readdata,
                                             nios_system_clock_10_in_waitrequest,
                                             reset_n,

                                            // outputs:
                                             cpu_2_data_master_byteenable_nios_system_clock_10_in,
                                             cpu_2_data_master_granted_nios_system_clock_10_in,
                                             cpu_2_data_master_qualified_request_nios_system_clock_10_in,
                                             cpu_2_data_master_read_data_valid_nios_system_clock_10_in,
                                             cpu_2_data_master_requests_nios_system_clock_10_in,
                                             d1_nios_system_clock_10_in_end_xfer,
                                             nios_system_clock_10_in_address,
                                             nios_system_clock_10_in_endofpacket_from_sa,
                                             nios_system_clock_10_in_nativeaddress,
                                             nios_system_clock_10_in_read,
                                             nios_system_clock_10_in_readdata_from_sa,
                                             nios_system_clock_10_in_reset_n,
                                             nios_system_clock_10_in_waitrequest_from_sa,
                                             nios_system_clock_10_in_write,
                                             nios_system_clock_10_in_writedata
                                          )
;

  output           cpu_2_data_master_byteenable_nios_system_clock_10_in;
  output           cpu_2_data_master_granted_nios_system_clock_10_in;
  output           cpu_2_data_master_qualified_request_nios_system_clock_10_in;
  output           cpu_2_data_master_read_data_valid_nios_system_clock_10_in;
  output           cpu_2_data_master_requests_nios_system_clock_10_in;
  output           d1_nios_system_clock_10_in_end_xfer;
  output           nios_system_clock_10_in_address;
  output           nios_system_clock_10_in_endofpacket_from_sa;
  output           nios_system_clock_10_in_nativeaddress;
  output           nios_system_clock_10_in_read;
  output  [  7: 0] nios_system_clock_10_in_readdata_from_sa;
  output           nios_system_clock_10_in_reset_n;
  output           nios_system_clock_10_in_waitrequest_from_sa;
  output           nios_system_clock_10_in_write;
  output  [  7: 0] nios_system_clock_10_in_writedata;
  input            clk;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input   [  3: 0] cpu_2_data_master_byteenable;
  input   [  1: 0] cpu_2_data_master_dbs_address;
  input   [  7: 0] cpu_2_data_master_dbs_write_8;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input            nios_system_clock_10_in_endofpacket;
  input   [  7: 0] nios_system_clock_10_in_readdata;
  input            nios_system_clock_10_in_waitrequest;
  input            reset_n;

  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_byteenable_nios_system_clock_10_in;
  wire             cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_0;
  wire             cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_1;
  wire             cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_2;
  wire             cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_3;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_nios_system_clock_10_in;
  wire             cpu_2_data_master_qualified_request_nios_system_clock_10_in;
  wire             cpu_2_data_master_read_data_valid_nios_system_clock_10_in;
  wire             cpu_2_data_master_requests_nios_system_clock_10_in;
  wire             cpu_2_data_master_saved_grant_nios_system_clock_10_in;
  reg              d1_nios_system_clock_10_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_10_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             nios_system_clock_10_in_address;
  wire             nios_system_clock_10_in_allgrants;
  wire             nios_system_clock_10_in_allow_new_arb_cycle;
  wire             nios_system_clock_10_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_10_in_any_continuerequest;
  wire             nios_system_clock_10_in_arb_counter_enable;
  reg     [  2: 0] nios_system_clock_10_in_arb_share_counter;
  wire    [  2: 0] nios_system_clock_10_in_arb_share_counter_next_value;
  wire    [  2: 0] nios_system_clock_10_in_arb_share_set_values;
  wire             nios_system_clock_10_in_beginbursttransfer_internal;
  wire             nios_system_clock_10_in_begins_xfer;
  wire             nios_system_clock_10_in_end_xfer;
  wire             nios_system_clock_10_in_endofpacket_from_sa;
  wire             nios_system_clock_10_in_firsttransfer;
  wire             nios_system_clock_10_in_grant_vector;
  wire             nios_system_clock_10_in_in_a_read_cycle;
  wire             nios_system_clock_10_in_in_a_write_cycle;
  wire             nios_system_clock_10_in_master_qreq_vector;
  wire             nios_system_clock_10_in_nativeaddress;
  wire             nios_system_clock_10_in_non_bursting_master_requests;
  wire             nios_system_clock_10_in_pretend_byte_enable;
  wire             nios_system_clock_10_in_read;
  wire    [  7: 0] nios_system_clock_10_in_readdata_from_sa;
  reg              nios_system_clock_10_in_reg_firsttransfer;
  wire             nios_system_clock_10_in_reset_n;
  reg              nios_system_clock_10_in_slavearbiterlockenable;
  wire             nios_system_clock_10_in_slavearbiterlockenable2;
  wire             nios_system_clock_10_in_unreg_firsttransfer;
  wire             nios_system_clock_10_in_waitrequest_from_sa;
  wire             nios_system_clock_10_in_waits_for_read;
  wire             nios_system_clock_10_in_waits_for_write;
  wire             nios_system_clock_10_in_write;
  wire    [  7: 0] nios_system_clock_10_in_writedata;
  wire             wait_for_nios_system_clock_10_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_10_in_end_xfer;
    end


  assign nios_system_clock_10_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_2_data_master_qualified_request_nios_system_clock_10_in));
  //assign nios_system_clock_10_in_readdata_from_sa = nios_system_clock_10_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_10_in_readdata_from_sa = nios_system_clock_10_in_readdata;

  assign cpu_2_data_master_requests_nios_system_clock_10_in = ({cpu_2_data_master_address_to_slave[24 : 1] , 1'b0} == 25'h19030d8) & (cpu_2_data_master_read | cpu_2_data_master_write);
  //assign nios_system_clock_10_in_waitrequest_from_sa = nios_system_clock_10_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_10_in_waitrequest_from_sa = nios_system_clock_10_in_waitrequest;

  //nios_system_clock_10_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_10_in_arb_share_set_values = (cpu_2_data_master_granted_nios_system_clock_10_in)? 4 :
    1;

  //nios_system_clock_10_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_10_in_non_bursting_master_requests = cpu_2_data_master_requests_nios_system_clock_10_in;

  //nios_system_clock_10_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_10_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_10_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_10_in_arb_share_counter_next_value = nios_system_clock_10_in_firsttransfer ? (nios_system_clock_10_in_arb_share_set_values - 1) : |nios_system_clock_10_in_arb_share_counter ? (nios_system_clock_10_in_arb_share_counter - 1) : 0;

  //nios_system_clock_10_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_10_in_allgrants = |nios_system_clock_10_in_grant_vector;

  //nios_system_clock_10_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_10_in_end_xfer = ~(nios_system_clock_10_in_waits_for_read | nios_system_clock_10_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_10_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_10_in = nios_system_clock_10_in_end_xfer & (~nios_system_clock_10_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_10_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_10_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_10_in & nios_system_clock_10_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_10_in & ~nios_system_clock_10_in_non_bursting_master_requests);

  //nios_system_clock_10_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_10_in_arb_share_counter <= 0;
      else if (nios_system_clock_10_in_arb_counter_enable)
          nios_system_clock_10_in_arb_share_counter <= nios_system_clock_10_in_arb_share_counter_next_value;
    end


  //nios_system_clock_10_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_10_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_10_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_10_in) | (end_xfer_arb_share_counter_term_nios_system_clock_10_in & ~nios_system_clock_10_in_non_bursting_master_requests))
          nios_system_clock_10_in_slavearbiterlockenable <= |nios_system_clock_10_in_arb_share_counter_next_value;
    end


  //cpu_2/data_master nios_system_clock_10/in arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = nios_system_clock_10_in_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //nios_system_clock_10_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_10_in_slavearbiterlockenable2 = |nios_system_clock_10_in_arb_share_counter_next_value;

  //cpu_2/data_master nios_system_clock_10/in arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = nios_system_clock_10_in_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //nios_system_clock_10_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_10_in_any_continuerequest = 1;

  //cpu_2_data_master_continuerequest continued request, which is an e_assign
  assign cpu_2_data_master_continuerequest = 1;

  assign cpu_2_data_master_qualified_request_nios_system_clock_10_in = cpu_2_data_master_requests_nios_system_clock_10_in & ~((cpu_2_data_master_read & ((cpu_2_data_master_latency_counter != 0) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | ((!cpu_2_data_master_byteenable_nios_system_clock_10_in) & cpu_2_data_master_write));
  //local readdatavalid cpu_2_data_master_read_data_valid_nios_system_clock_10_in, which is an e_mux
  assign cpu_2_data_master_read_data_valid_nios_system_clock_10_in = cpu_2_data_master_granted_nios_system_clock_10_in & cpu_2_data_master_read & ~nios_system_clock_10_in_waits_for_read;

  //nios_system_clock_10_in_writedata mux, which is an e_mux
  assign nios_system_clock_10_in_writedata = cpu_2_data_master_dbs_write_8;

  //assign nios_system_clock_10_in_endofpacket_from_sa = nios_system_clock_10_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_10_in_endofpacket_from_sa = nios_system_clock_10_in_endofpacket;

  //master is always granted when requested
  assign cpu_2_data_master_granted_nios_system_clock_10_in = cpu_2_data_master_qualified_request_nios_system_clock_10_in;

  //cpu_2/data_master saved-grant nios_system_clock_10/in, which is an e_assign
  assign cpu_2_data_master_saved_grant_nios_system_clock_10_in = cpu_2_data_master_requests_nios_system_clock_10_in;

  //allow new arb cycle for nios_system_clock_10/in, which is an e_assign
  assign nios_system_clock_10_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_10_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_10_in_master_qreq_vector = 1;

  //nios_system_clock_10_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_10_in_reset_n = reset_n;

  //nios_system_clock_10_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_10_in_firsttransfer = nios_system_clock_10_in_begins_xfer ? nios_system_clock_10_in_unreg_firsttransfer : nios_system_clock_10_in_reg_firsttransfer;

  //nios_system_clock_10_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_10_in_unreg_firsttransfer = ~(nios_system_clock_10_in_slavearbiterlockenable & nios_system_clock_10_in_any_continuerequest);

  //nios_system_clock_10_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_10_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_10_in_begins_xfer)
          nios_system_clock_10_in_reg_firsttransfer <= nios_system_clock_10_in_unreg_firsttransfer;
    end


  //nios_system_clock_10_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_10_in_beginbursttransfer_internal = nios_system_clock_10_in_begins_xfer;

  //nios_system_clock_10_in_read assignment, which is an e_mux
  assign nios_system_clock_10_in_read = cpu_2_data_master_granted_nios_system_clock_10_in & cpu_2_data_master_read;

  //nios_system_clock_10_in_write assignment, which is an e_mux
  assign nios_system_clock_10_in_write = ((cpu_2_data_master_granted_nios_system_clock_10_in & cpu_2_data_master_write)) & nios_system_clock_10_in_pretend_byte_enable;

  //nios_system_clock_10_in_address mux, which is an e_mux
  assign nios_system_clock_10_in_address = {cpu_2_data_master_address_to_slave >> 2,
    cpu_2_data_master_dbs_address[1 : 0]};

  //slaveid nios_system_clock_10_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_10_in_nativeaddress = cpu_2_data_master_address_to_slave >> 2;

  //d1_nios_system_clock_10_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_10_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_10_in_end_xfer <= nios_system_clock_10_in_end_xfer;
    end


  //nios_system_clock_10_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_10_in_waits_for_read = nios_system_clock_10_in_in_a_read_cycle & nios_system_clock_10_in_waitrequest_from_sa;

  //nios_system_clock_10_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_10_in_in_a_read_cycle = cpu_2_data_master_granted_nios_system_clock_10_in & cpu_2_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_10_in_in_a_read_cycle;

  //nios_system_clock_10_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_10_in_waits_for_write = nios_system_clock_10_in_in_a_write_cycle & nios_system_clock_10_in_waitrequest_from_sa;

  //nios_system_clock_10_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_10_in_in_a_write_cycle = cpu_2_data_master_granted_nios_system_clock_10_in & cpu_2_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_10_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_10_in_counter = 0;
  //nios_system_clock_10_in_pretend_byte_enable byte enable port mux, which is an e_mux
  assign nios_system_clock_10_in_pretend_byte_enable = (cpu_2_data_master_granted_nios_system_clock_10_in)? cpu_2_data_master_byteenable_nios_system_clock_10_in :
    -1;

  assign {cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_3,
cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_2,
cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_1,
cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_0} = cpu_2_data_master_byteenable;
  assign cpu_2_data_master_byteenable_nios_system_clock_10_in = ((cpu_2_data_master_dbs_address[1 : 0] == 0))? cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_0 :
    ((cpu_2_data_master_dbs_address[1 : 0] == 1))? cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_1 :
    ((cpu_2_data_master_dbs_address[1 : 0] == 2))? cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_2 :
    cpu_2_data_master_byteenable_nios_system_clock_10_in_segment_3;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_10/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_10_out_arbitrator (
                                             // inputs:
                                              clk,
                                              clocks_0_avalon_clocks_slave_readdata_from_sa,
                                              d1_clocks_0_avalon_clocks_slave_end_xfer,
                                              nios_system_clock_10_out_address,
                                              nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave,
                                              nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave,
                                              nios_system_clock_10_out_read,
                                              nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave,
                                              nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave,
                                              nios_system_clock_10_out_write,
                                              nios_system_clock_10_out_writedata,
                                              reset_n,

                                             // outputs:
                                              nios_system_clock_10_out_address_to_slave,
                                              nios_system_clock_10_out_readdata,
                                              nios_system_clock_10_out_reset_n,
                                              nios_system_clock_10_out_waitrequest
                                           )
;

  output           nios_system_clock_10_out_address_to_slave;
  output  [  7: 0] nios_system_clock_10_out_readdata;
  output           nios_system_clock_10_out_reset_n;
  output           nios_system_clock_10_out_waitrequest;
  input            clk;
  input   [  7: 0] clocks_0_avalon_clocks_slave_readdata_from_sa;
  input            d1_clocks_0_avalon_clocks_slave_end_xfer;
  input            nios_system_clock_10_out_address;
  input            nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_10_out_read;
  input            nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_10_out_write;
  input   [  7: 0] nios_system_clock_10_out_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg              nios_system_clock_10_out_address_last_time;
  wire             nios_system_clock_10_out_address_to_slave;
  reg              nios_system_clock_10_out_read_last_time;
  wire    [  7: 0] nios_system_clock_10_out_readdata;
  wire             nios_system_clock_10_out_reset_n;
  wire             nios_system_clock_10_out_run;
  wire             nios_system_clock_10_out_waitrequest;
  reg              nios_system_clock_10_out_write_last_time;
  reg     [  7: 0] nios_system_clock_10_out_writedata_last_time;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave | nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave | ~nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave) & (nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave | ~nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave) & ((~nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave | ~nios_system_clock_10_out_read | (nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave & nios_system_clock_10_out_read))) & ((~nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave | ~(nios_system_clock_10_out_read | nios_system_clock_10_out_write) | (1 & (nios_system_clock_10_out_read | nios_system_clock_10_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_10_out_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_10_out_address_to_slave = nios_system_clock_10_out_address;

  //nios_system_clock_10/out readdata mux, which is an e_mux
  assign nios_system_clock_10_out_readdata = clocks_0_avalon_clocks_slave_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_10_out_waitrequest = ~nios_system_clock_10_out_run;

  //nios_system_clock_10_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_10_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_10_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_10_out_address_last_time <= 0;
      else 
        nios_system_clock_10_out_address_last_time <= nios_system_clock_10_out_address;
    end


  //nios_system_clock_10/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_10_out_waitrequest & (nios_system_clock_10_out_read | nios_system_clock_10_out_write);
    end


  //nios_system_clock_10_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_10_out_address != nios_system_clock_10_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_10_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_10_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_10_out_read_last_time <= 0;
      else 
        nios_system_clock_10_out_read_last_time <= nios_system_clock_10_out_read;
    end


  //nios_system_clock_10_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_10_out_read != nios_system_clock_10_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_10_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_10_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_10_out_write_last_time <= 0;
      else 
        nios_system_clock_10_out_write_last_time <= nios_system_clock_10_out_write;
    end


  //nios_system_clock_10_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_10_out_write != nios_system_clock_10_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_10_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_10_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_10_out_writedata_last_time <= 0;
      else 
        nios_system_clock_10_out_writedata_last_time <= nios_system_clock_10_out_writedata;
    end


  //nios_system_clock_10_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_10_out_writedata != nios_system_clock_10_out_writedata_last_time) & nios_system_clock_10_out_write)
        begin
          $write("%0d ns: nios_system_clock_10_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_11_in_arbitrator (
                                            // inputs:
                                             clk,
                                             cpu_3_data_master_address_to_slave,
                                             cpu_3_data_master_byteenable,
                                             cpu_3_data_master_dbs_address,
                                             cpu_3_data_master_dbs_write_8,
                                             cpu_3_data_master_latency_counter,
                                             cpu_3_data_master_read,
                                             cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                             cpu_3_data_master_write,
                                             nios_system_clock_11_in_endofpacket,
                                             nios_system_clock_11_in_readdata,
                                             nios_system_clock_11_in_waitrequest,
                                             reset_n,

                                            // outputs:
                                             cpu_3_data_master_byteenable_nios_system_clock_11_in,
                                             cpu_3_data_master_granted_nios_system_clock_11_in,
                                             cpu_3_data_master_qualified_request_nios_system_clock_11_in,
                                             cpu_3_data_master_read_data_valid_nios_system_clock_11_in,
                                             cpu_3_data_master_requests_nios_system_clock_11_in,
                                             d1_nios_system_clock_11_in_end_xfer,
                                             nios_system_clock_11_in_address,
                                             nios_system_clock_11_in_endofpacket_from_sa,
                                             nios_system_clock_11_in_nativeaddress,
                                             nios_system_clock_11_in_read,
                                             nios_system_clock_11_in_readdata_from_sa,
                                             nios_system_clock_11_in_reset_n,
                                             nios_system_clock_11_in_waitrequest_from_sa,
                                             nios_system_clock_11_in_write,
                                             nios_system_clock_11_in_writedata
                                          )
;

  output           cpu_3_data_master_byteenable_nios_system_clock_11_in;
  output           cpu_3_data_master_granted_nios_system_clock_11_in;
  output           cpu_3_data_master_qualified_request_nios_system_clock_11_in;
  output           cpu_3_data_master_read_data_valid_nios_system_clock_11_in;
  output           cpu_3_data_master_requests_nios_system_clock_11_in;
  output           d1_nios_system_clock_11_in_end_xfer;
  output           nios_system_clock_11_in_address;
  output           nios_system_clock_11_in_endofpacket_from_sa;
  output           nios_system_clock_11_in_nativeaddress;
  output           nios_system_clock_11_in_read;
  output  [  7: 0] nios_system_clock_11_in_readdata_from_sa;
  output           nios_system_clock_11_in_reset_n;
  output           nios_system_clock_11_in_waitrequest_from_sa;
  output           nios_system_clock_11_in_write;
  output  [  7: 0] nios_system_clock_11_in_writedata;
  input            clk;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input   [  3: 0] cpu_3_data_master_byteenable;
  input   [  1: 0] cpu_3_data_master_dbs_address;
  input   [  7: 0] cpu_3_data_master_dbs_write_8;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input            nios_system_clock_11_in_endofpacket;
  input   [  7: 0] nios_system_clock_11_in_readdata;
  input            nios_system_clock_11_in_waitrequest;
  input            reset_n;

  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_byteenable_nios_system_clock_11_in;
  wire             cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_0;
  wire             cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_1;
  wire             cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_2;
  wire             cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_3;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_nios_system_clock_11_in;
  wire             cpu_3_data_master_qualified_request_nios_system_clock_11_in;
  wire             cpu_3_data_master_read_data_valid_nios_system_clock_11_in;
  wire             cpu_3_data_master_requests_nios_system_clock_11_in;
  wire             cpu_3_data_master_saved_grant_nios_system_clock_11_in;
  reg              d1_nios_system_clock_11_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_11_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             nios_system_clock_11_in_address;
  wire             nios_system_clock_11_in_allgrants;
  wire             nios_system_clock_11_in_allow_new_arb_cycle;
  wire             nios_system_clock_11_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_11_in_any_continuerequest;
  wire             nios_system_clock_11_in_arb_counter_enable;
  reg     [  2: 0] nios_system_clock_11_in_arb_share_counter;
  wire    [  2: 0] nios_system_clock_11_in_arb_share_counter_next_value;
  wire    [  2: 0] nios_system_clock_11_in_arb_share_set_values;
  wire             nios_system_clock_11_in_beginbursttransfer_internal;
  wire             nios_system_clock_11_in_begins_xfer;
  wire             nios_system_clock_11_in_end_xfer;
  wire             nios_system_clock_11_in_endofpacket_from_sa;
  wire             nios_system_clock_11_in_firsttransfer;
  wire             nios_system_clock_11_in_grant_vector;
  wire             nios_system_clock_11_in_in_a_read_cycle;
  wire             nios_system_clock_11_in_in_a_write_cycle;
  wire             nios_system_clock_11_in_master_qreq_vector;
  wire             nios_system_clock_11_in_nativeaddress;
  wire             nios_system_clock_11_in_non_bursting_master_requests;
  wire             nios_system_clock_11_in_pretend_byte_enable;
  wire             nios_system_clock_11_in_read;
  wire    [  7: 0] nios_system_clock_11_in_readdata_from_sa;
  reg              nios_system_clock_11_in_reg_firsttransfer;
  wire             nios_system_clock_11_in_reset_n;
  reg              nios_system_clock_11_in_slavearbiterlockenable;
  wire             nios_system_clock_11_in_slavearbiterlockenable2;
  wire             nios_system_clock_11_in_unreg_firsttransfer;
  wire             nios_system_clock_11_in_waitrequest_from_sa;
  wire             nios_system_clock_11_in_waits_for_read;
  wire             nios_system_clock_11_in_waits_for_write;
  wire             nios_system_clock_11_in_write;
  wire    [  7: 0] nios_system_clock_11_in_writedata;
  wire             wait_for_nios_system_clock_11_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_11_in_end_xfer;
    end


  assign nios_system_clock_11_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_3_data_master_qualified_request_nios_system_clock_11_in));
  //assign nios_system_clock_11_in_readdata_from_sa = nios_system_clock_11_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_11_in_readdata_from_sa = nios_system_clock_11_in_readdata;

  assign cpu_3_data_master_requests_nios_system_clock_11_in = ({cpu_3_data_master_address_to_slave[24 : 1] , 1'b0} == 25'h19030d8) & (cpu_3_data_master_read | cpu_3_data_master_write);
  //assign nios_system_clock_11_in_waitrequest_from_sa = nios_system_clock_11_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_11_in_waitrequest_from_sa = nios_system_clock_11_in_waitrequest;

  //nios_system_clock_11_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_11_in_arb_share_set_values = (cpu_3_data_master_granted_nios_system_clock_11_in)? 4 :
    1;

  //nios_system_clock_11_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_11_in_non_bursting_master_requests = cpu_3_data_master_requests_nios_system_clock_11_in;

  //nios_system_clock_11_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_11_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_11_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_11_in_arb_share_counter_next_value = nios_system_clock_11_in_firsttransfer ? (nios_system_clock_11_in_arb_share_set_values - 1) : |nios_system_clock_11_in_arb_share_counter ? (nios_system_clock_11_in_arb_share_counter - 1) : 0;

  //nios_system_clock_11_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_11_in_allgrants = |nios_system_clock_11_in_grant_vector;

  //nios_system_clock_11_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_11_in_end_xfer = ~(nios_system_clock_11_in_waits_for_read | nios_system_clock_11_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_11_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_11_in = nios_system_clock_11_in_end_xfer & (~nios_system_clock_11_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_11_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_11_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_11_in & nios_system_clock_11_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_11_in & ~nios_system_clock_11_in_non_bursting_master_requests);

  //nios_system_clock_11_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_11_in_arb_share_counter <= 0;
      else if (nios_system_clock_11_in_arb_counter_enable)
          nios_system_clock_11_in_arb_share_counter <= nios_system_clock_11_in_arb_share_counter_next_value;
    end


  //nios_system_clock_11_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_11_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_11_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_11_in) | (end_xfer_arb_share_counter_term_nios_system_clock_11_in & ~nios_system_clock_11_in_non_bursting_master_requests))
          nios_system_clock_11_in_slavearbiterlockenable <= |nios_system_clock_11_in_arb_share_counter_next_value;
    end


  //cpu_3/data_master nios_system_clock_11/in arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = nios_system_clock_11_in_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //nios_system_clock_11_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_11_in_slavearbiterlockenable2 = |nios_system_clock_11_in_arb_share_counter_next_value;

  //cpu_3/data_master nios_system_clock_11/in arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = nios_system_clock_11_in_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //nios_system_clock_11_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_11_in_any_continuerequest = 1;

  //cpu_3_data_master_continuerequest continued request, which is an e_assign
  assign cpu_3_data_master_continuerequest = 1;

  assign cpu_3_data_master_qualified_request_nios_system_clock_11_in = cpu_3_data_master_requests_nios_system_clock_11_in & ~((cpu_3_data_master_read & ((cpu_3_data_master_latency_counter != 0) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | ((!cpu_3_data_master_byteenable_nios_system_clock_11_in) & cpu_3_data_master_write));
  //local readdatavalid cpu_3_data_master_read_data_valid_nios_system_clock_11_in, which is an e_mux
  assign cpu_3_data_master_read_data_valid_nios_system_clock_11_in = cpu_3_data_master_granted_nios_system_clock_11_in & cpu_3_data_master_read & ~nios_system_clock_11_in_waits_for_read;

  //nios_system_clock_11_in_writedata mux, which is an e_mux
  assign nios_system_clock_11_in_writedata = cpu_3_data_master_dbs_write_8;

  //assign nios_system_clock_11_in_endofpacket_from_sa = nios_system_clock_11_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_11_in_endofpacket_from_sa = nios_system_clock_11_in_endofpacket;

  //master is always granted when requested
  assign cpu_3_data_master_granted_nios_system_clock_11_in = cpu_3_data_master_qualified_request_nios_system_clock_11_in;

  //cpu_3/data_master saved-grant nios_system_clock_11/in, which is an e_assign
  assign cpu_3_data_master_saved_grant_nios_system_clock_11_in = cpu_3_data_master_requests_nios_system_clock_11_in;

  //allow new arb cycle for nios_system_clock_11/in, which is an e_assign
  assign nios_system_clock_11_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_11_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_11_in_master_qreq_vector = 1;

  //nios_system_clock_11_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_11_in_reset_n = reset_n;

  //nios_system_clock_11_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_11_in_firsttransfer = nios_system_clock_11_in_begins_xfer ? nios_system_clock_11_in_unreg_firsttransfer : nios_system_clock_11_in_reg_firsttransfer;

  //nios_system_clock_11_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_11_in_unreg_firsttransfer = ~(nios_system_clock_11_in_slavearbiterlockenable & nios_system_clock_11_in_any_continuerequest);

  //nios_system_clock_11_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_11_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_11_in_begins_xfer)
          nios_system_clock_11_in_reg_firsttransfer <= nios_system_clock_11_in_unreg_firsttransfer;
    end


  //nios_system_clock_11_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_11_in_beginbursttransfer_internal = nios_system_clock_11_in_begins_xfer;

  //nios_system_clock_11_in_read assignment, which is an e_mux
  assign nios_system_clock_11_in_read = cpu_3_data_master_granted_nios_system_clock_11_in & cpu_3_data_master_read;

  //nios_system_clock_11_in_write assignment, which is an e_mux
  assign nios_system_clock_11_in_write = ((cpu_3_data_master_granted_nios_system_clock_11_in & cpu_3_data_master_write)) & nios_system_clock_11_in_pretend_byte_enable;

  //nios_system_clock_11_in_address mux, which is an e_mux
  assign nios_system_clock_11_in_address = {cpu_3_data_master_address_to_slave >> 2,
    cpu_3_data_master_dbs_address[1 : 0]};

  //slaveid nios_system_clock_11_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_11_in_nativeaddress = cpu_3_data_master_address_to_slave >> 2;

  //d1_nios_system_clock_11_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_11_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_11_in_end_xfer <= nios_system_clock_11_in_end_xfer;
    end


  //nios_system_clock_11_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_11_in_waits_for_read = nios_system_clock_11_in_in_a_read_cycle & nios_system_clock_11_in_waitrequest_from_sa;

  //nios_system_clock_11_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_11_in_in_a_read_cycle = cpu_3_data_master_granted_nios_system_clock_11_in & cpu_3_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_11_in_in_a_read_cycle;

  //nios_system_clock_11_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_11_in_waits_for_write = nios_system_clock_11_in_in_a_write_cycle & nios_system_clock_11_in_waitrequest_from_sa;

  //nios_system_clock_11_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_11_in_in_a_write_cycle = cpu_3_data_master_granted_nios_system_clock_11_in & cpu_3_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_11_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_11_in_counter = 0;
  //nios_system_clock_11_in_pretend_byte_enable byte enable port mux, which is an e_mux
  assign nios_system_clock_11_in_pretend_byte_enable = (cpu_3_data_master_granted_nios_system_clock_11_in)? cpu_3_data_master_byteenable_nios_system_clock_11_in :
    -1;

  assign {cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_3,
cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_2,
cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_1,
cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_0} = cpu_3_data_master_byteenable;
  assign cpu_3_data_master_byteenable_nios_system_clock_11_in = ((cpu_3_data_master_dbs_address[1 : 0] == 0))? cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_0 :
    ((cpu_3_data_master_dbs_address[1 : 0] == 1))? cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_1 :
    ((cpu_3_data_master_dbs_address[1 : 0] == 2))? cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_2 :
    cpu_3_data_master_byteenable_nios_system_clock_11_in_segment_3;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_11/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_11_out_arbitrator (
                                             // inputs:
                                              clk,
                                              clocks_0_avalon_clocks_slave_readdata_from_sa,
                                              d1_clocks_0_avalon_clocks_slave_end_xfer,
                                              nios_system_clock_11_out_address,
                                              nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave,
                                              nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave,
                                              nios_system_clock_11_out_read,
                                              nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave,
                                              nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave,
                                              nios_system_clock_11_out_write,
                                              nios_system_clock_11_out_writedata,
                                              reset_n,

                                             // outputs:
                                              nios_system_clock_11_out_address_to_slave,
                                              nios_system_clock_11_out_readdata,
                                              nios_system_clock_11_out_reset_n,
                                              nios_system_clock_11_out_waitrequest
                                           )
;

  output           nios_system_clock_11_out_address_to_slave;
  output  [  7: 0] nios_system_clock_11_out_readdata;
  output           nios_system_clock_11_out_reset_n;
  output           nios_system_clock_11_out_waitrequest;
  input            clk;
  input   [  7: 0] clocks_0_avalon_clocks_slave_readdata_from_sa;
  input            d1_clocks_0_avalon_clocks_slave_end_xfer;
  input            nios_system_clock_11_out_address;
  input            nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_11_out_read;
  input            nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_11_out_write;
  input   [  7: 0] nios_system_clock_11_out_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg              nios_system_clock_11_out_address_last_time;
  wire             nios_system_clock_11_out_address_to_slave;
  reg              nios_system_clock_11_out_read_last_time;
  wire    [  7: 0] nios_system_clock_11_out_readdata;
  wire             nios_system_clock_11_out_reset_n;
  wire             nios_system_clock_11_out_run;
  wire             nios_system_clock_11_out_waitrequest;
  reg              nios_system_clock_11_out_write_last_time;
  reg     [  7: 0] nios_system_clock_11_out_writedata_last_time;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave | nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave | ~nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave) & (nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave | ~nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave) & ((~nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave | ~nios_system_clock_11_out_read | (nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave & nios_system_clock_11_out_read))) & ((~nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave | ~(nios_system_clock_11_out_read | nios_system_clock_11_out_write) | (1 & (nios_system_clock_11_out_read | nios_system_clock_11_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_11_out_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_11_out_address_to_slave = nios_system_clock_11_out_address;

  //nios_system_clock_11/out readdata mux, which is an e_mux
  assign nios_system_clock_11_out_readdata = clocks_0_avalon_clocks_slave_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_11_out_waitrequest = ~nios_system_clock_11_out_run;

  //nios_system_clock_11_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_11_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_11_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_11_out_address_last_time <= 0;
      else 
        nios_system_clock_11_out_address_last_time <= nios_system_clock_11_out_address;
    end


  //nios_system_clock_11/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_11_out_waitrequest & (nios_system_clock_11_out_read | nios_system_clock_11_out_write);
    end


  //nios_system_clock_11_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_11_out_address != nios_system_clock_11_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_11_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_11_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_11_out_read_last_time <= 0;
      else 
        nios_system_clock_11_out_read_last_time <= nios_system_clock_11_out_read;
    end


  //nios_system_clock_11_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_11_out_read != nios_system_clock_11_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_11_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_11_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_11_out_write_last_time <= 0;
      else 
        nios_system_clock_11_out_write_last_time <= nios_system_clock_11_out_write;
    end


  //nios_system_clock_11_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_11_out_write != nios_system_clock_11_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_11_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_11_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_11_out_writedata_last_time <= 0;
      else 
        nios_system_clock_11_out_writedata_last_time <= nios_system_clock_11_out_writedata;
    end


  //nios_system_clock_11_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_11_out_writedata != nios_system_clock_11_out_writedata_last_time) & nios_system_clock_11_out_write)
        begin
          $write("%0d ns: nios_system_clock_11_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_2_in_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_0_instruction_master_address_to_slave,
                                            cpu_0_instruction_master_dbs_address,
                                            cpu_0_instruction_master_latency_counter,
                                            cpu_0_instruction_master_read,
                                            nios_system_clock_2_in_endofpacket,
                                            nios_system_clock_2_in_readdata,
                                            nios_system_clock_2_in_waitrequest,
                                            reset_n,

                                           // outputs:
                                            cpu_0_instruction_master_granted_nios_system_clock_2_in,
                                            cpu_0_instruction_master_qualified_request_nios_system_clock_2_in,
                                            cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in,
                                            cpu_0_instruction_master_requests_nios_system_clock_2_in,
                                            d1_nios_system_clock_2_in_end_xfer,
                                            nios_system_clock_2_in_address,
                                            nios_system_clock_2_in_byteenable,
                                            nios_system_clock_2_in_endofpacket_from_sa,
                                            nios_system_clock_2_in_nativeaddress,
                                            nios_system_clock_2_in_read,
                                            nios_system_clock_2_in_readdata_from_sa,
                                            nios_system_clock_2_in_reset_n,
                                            nios_system_clock_2_in_waitrequest_from_sa,
                                            nios_system_clock_2_in_write
                                         )
;

  output           cpu_0_instruction_master_granted_nios_system_clock_2_in;
  output           cpu_0_instruction_master_qualified_request_nios_system_clock_2_in;
  output           cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in;
  output           cpu_0_instruction_master_requests_nios_system_clock_2_in;
  output           d1_nios_system_clock_2_in_end_xfer;
  output  [ 22: 0] nios_system_clock_2_in_address;
  output  [  1: 0] nios_system_clock_2_in_byteenable;
  output           nios_system_clock_2_in_endofpacket_from_sa;
  output  [ 21: 0] nios_system_clock_2_in_nativeaddress;
  output           nios_system_clock_2_in_read;
  output  [ 15: 0] nios_system_clock_2_in_readdata_from_sa;
  output           nios_system_clock_2_in_reset_n;
  output           nios_system_clock_2_in_waitrequest_from_sa;
  output           nios_system_clock_2_in_write;
  input            clk;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input   [  1: 0] cpu_0_instruction_master_dbs_address;
  input            cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input            nios_system_clock_2_in_endofpacket;
  input   [ 15: 0] nios_system_clock_2_in_readdata;
  input            nios_system_clock_2_in_waitrequest;
  input            reset_n;

  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_nios_system_clock_2_in;
  wire             cpu_0_instruction_master_qualified_request_nios_system_clock_2_in;
  wire             cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in;
  wire             cpu_0_instruction_master_requests_nios_system_clock_2_in;
  wire             cpu_0_instruction_master_saved_grant_nios_system_clock_2_in;
  reg              d1_nios_system_clock_2_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_2_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 22: 0] nios_system_clock_2_in_address;
  wire             nios_system_clock_2_in_allgrants;
  wire             nios_system_clock_2_in_allow_new_arb_cycle;
  wire             nios_system_clock_2_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_2_in_any_continuerequest;
  wire             nios_system_clock_2_in_arb_counter_enable;
  reg     [  1: 0] nios_system_clock_2_in_arb_share_counter;
  wire    [  1: 0] nios_system_clock_2_in_arb_share_counter_next_value;
  wire    [  1: 0] nios_system_clock_2_in_arb_share_set_values;
  wire             nios_system_clock_2_in_beginbursttransfer_internal;
  wire             nios_system_clock_2_in_begins_xfer;
  wire    [  1: 0] nios_system_clock_2_in_byteenable;
  wire             nios_system_clock_2_in_end_xfer;
  wire             nios_system_clock_2_in_endofpacket_from_sa;
  wire             nios_system_clock_2_in_firsttransfer;
  wire             nios_system_clock_2_in_grant_vector;
  wire             nios_system_clock_2_in_in_a_read_cycle;
  wire             nios_system_clock_2_in_in_a_write_cycle;
  wire             nios_system_clock_2_in_master_qreq_vector;
  wire    [ 21: 0] nios_system_clock_2_in_nativeaddress;
  wire             nios_system_clock_2_in_non_bursting_master_requests;
  wire             nios_system_clock_2_in_read;
  wire    [ 15: 0] nios_system_clock_2_in_readdata_from_sa;
  reg              nios_system_clock_2_in_reg_firsttransfer;
  wire             nios_system_clock_2_in_reset_n;
  reg              nios_system_clock_2_in_slavearbiterlockenable;
  wire             nios_system_clock_2_in_slavearbiterlockenable2;
  wire             nios_system_clock_2_in_unreg_firsttransfer;
  wire             nios_system_clock_2_in_waitrequest_from_sa;
  wire             nios_system_clock_2_in_waits_for_read;
  wire             nios_system_clock_2_in_waits_for_write;
  wire             nios_system_clock_2_in_write;
  wire             wait_for_nios_system_clock_2_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_2_in_end_xfer;
    end


  assign nios_system_clock_2_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_instruction_master_qualified_request_nios_system_clock_2_in));
  //assign nios_system_clock_2_in_readdata_from_sa = nios_system_clock_2_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_2_in_readdata_from_sa = nios_system_clock_2_in_readdata;

  assign cpu_0_instruction_master_requests_nios_system_clock_2_in = (({cpu_0_instruction_master_address_to_slave[24 : 23] , 23'b0} == 25'h800000) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //assign nios_system_clock_2_in_waitrequest_from_sa = nios_system_clock_2_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_2_in_waitrequest_from_sa = nios_system_clock_2_in_waitrequest;

  //nios_system_clock_2_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_2_in_arb_share_set_values = (cpu_0_instruction_master_granted_nios_system_clock_2_in)? 2 :
    1;

  //nios_system_clock_2_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_2_in_non_bursting_master_requests = cpu_0_instruction_master_requests_nios_system_clock_2_in;

  //nios_system_clock_2_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_2_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_2_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_2_in_arb_share_counter_next_value = nios_system_clock_2_in_firsttransfer ? (nios_system_clock_2_in_arb_share_set_values - 1) : |nios_system_clock_2_in_arb_share_counter ? (nios_system_clock_2_in_arb_share_counter - 1) : 0;

  //nios_system_clock_2_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_2_in_allgrants = |nios_system_clock_2_in_grant_vector;

  //nios_system_clock_2_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_2_in_end_xfer = ~(nios_system_clock_2_in_waits_for_read | nios_system_clock_2_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_2_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_2_in = nios_system_clock_2_in_end_xfer & (~nios_system_clock_2_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_2_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_2_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_2_in & nios_system_clock_2_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_2_in & ~nios_system_clock_2_in_non_bursting_master_requests);

  //nios_system_clock_2_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_2_in_arb_share_counter <= 0;
      else if (nios_system_clock_2_in_arb_counter_enable)
          nios_system_clock_2_in_arb_share_counter <= nios_system_clock_2_in_arb_share_counter_next_value;
    end


  //nios_system_clock_2_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_2_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_2_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_2_in) | (end_xfer_arb_share_counter_term_nios_system_clock_2_in & ~nios_system_clock_2_in_non_bursting_master_requests))
          nios_system_clock_2_in_slavearbiterlockenable <= |nios_system_clock_2_in_arb_share_counter_next_value;
    end


  //cpu_0/instruction_master nios_system_clock_2/in arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = nios_system_clock_2_in_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //nios_system_clock_2_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_2_in_slavearbiterlockenable2 = |nios_system_clock_2_in_arb_share_counter_next_value;

  //cpu_0/instruction_master nios_system_clock_2/in arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = nios_system_clock_2_in_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //nios_system_clock_2_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_2_in_any_continuerequest = 1;

  //cpu_0_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_0_instruction_master_continuerequest = 1;

  assign cpu_0_instruction_master_qualified_request_nios_system_clock_2_in = cpu_0_instruction_master_requests_nios_system_clock_2_in & ~((cpu_0_instruction_master_read & ((cpu_0_instruction_master_latency_counter != 0))));
  //local readdatavalid cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in = cpu_0_instruction_master_granted_nios_system_clock_2_in & cpu_0_instruction_master_read & ~nios_system_clock_2_in_waits_for_read;

  //assign nios_system_clock_2_in_endofpacket_from_sa = nios_system_clock_2_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_2_in_endofpacket_from_sa = nios_system_clock_2_in_endofpacket;

  //master is always granted when requested
  assign cpu_0_instruction_master_granted_nios_system_clock_2_in = cpu_0_instruction_master_qualified_request_nios_system_clock_2_in;

  //cpu_0/instruction_master saved-grant nios_system_clock_2/in, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_nios_system_clock_2_in = cpu_0_instruction_master_requests_nios_system_clock_2_in;

  //allow new arb cycle for nios_system_clock_2/in, which is an e_assign
  assign nios_system_clock_2_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_2_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_2_in_master_qreq_vector = 1;

  //nios_system_clock_2_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_2_in_reset_n = reset_n;

  //nios_system_clock_2_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_2_in_firsttransfer = nios_system_clock_2_in_begins_xfer ? nios_system_clock_2_in_unreg_firsttransfer : nios_system_clock_2_in_reg_firsttransfer;

  //nios_system_clock_2_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_2_in_unreg_firsttransfer = ~(nios_system_clock_2_in_slavearbiterlockenable & nios_system_clock_2_in_any_continuerequest);

  //nios_system_clock_2_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_2_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_2_in_begins_xfer)
          nios_system_clock_2_in_reg_firsttransfer <= nios_system_clock_2_in_unreg_firsttransfer;
    end


  //nios_system_clock_2_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_2_in_beginbursttransfer_internal = nios_system_clock_2_in_begins_xfer;

  //nios_system_clock_2_in_read assignment, which is an e_mux
  assign nios_system_clock_2_in_read = cpu_0_instruction_master_granted_nios_system_clock_2_in & cpu_0_instruction_master_read;

  //nios_system_clock_2_in_write assignment, which is an e_mux
  assign nios_system_clock_2_in_write = 0;

  //nios_system_clock_2_in_address mux, which is an e_mux
  assign nios_system_clock_2_in_address = {cpu_0_instruction_master_address_to_slave >> 2,
    cpu_0_instruction_master_dbs_address[1],
    {1 {1'b0}}};

  //slaveid nios_system_clock_2_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_2_in_nativeaddress = cpu_0_instruction_master_address_to_slave >> 2;

  //d1_nios_system_clock_2_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_2_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_2_in_end_xfer <= nios_system_clock_2_in_end_xfer;
    end


  //nios_system_clock_2_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_2_in_waits_for_read = nios_system_clock_2_in_in_a_read_cycle & nios_system_clock_2_in_waitrequest_from_sa;

  //nios_system_clock_2_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_2_in_in_a_read_cycle = cpu_0_instruction_master_granted_nios_system_clock_2_in & cpu_0_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_2_in_in_a_read_cycle;

  //nios_system_clock_2_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_2_in_waits_for_write = nios_system_clock_2_in_in_a_write_cycle & nios_system_clock_2_in_waitrequest_from_sa;

  //nios_system_clock_2_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_2_in_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_2_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_2_in_counter = 0;
  //nios_system_clock_2_in_byteenable byte enable port mux, which is an e_mux
  assign nios_system_clock_2_in_byteenable = -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_2/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_2_out_arbitrator (
                                            // inputs:
                                             clk,
                                             d1_sdram_0_s1_end_xfer,
                                             nios_system_clock_2_out_address,
                                             nios_system_clock_2_out_byteenable,
                                             nios_system_clock_2_out_granted_sdram_0_s1,
                                             nios_system_clock_2_out_qualified_request_sdram_0_s1,
                                             nios_system_clock_2_out_read,
                                             nios_system_clock_2_out_read_data_valid_sdram_0_s1,
                                             nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register,
                                             nios_system_clock_2_out_requests_sdram_0_s1,
                                             nios_system_clock_2_out_write,
                                             nios_system_clock_2_out_writedata,
                                             reset_n,
                                             sdram_0_s1_readdata_from_sa,
                                             sdram_0_s1_waitrequest_from_sa,

                                            // outputs:
                                             nios_system_clock_2_out_address_to_slave,
                                             nios_system_clock_2_out_readdata,
                                             nios_system_clock_2_out_reset_n,
                                             nios_system_clock_2_out_waitrequest
                                          )
;

  output  [ 22: 0] nios_system_clock_2_out_address_to_slave;
  output  [ 15: 0] nios_system_clock_2_out_readdata;
  output           nios_system_clock_2_out_reset_n;
  output           nios_system_clock_2_out_waitrequest;
  input            clk;
  input            d1_sdram_0_s1_end_xfer;
  input   [ 22: 0] nios_system_clock_2_out_address;
  input   [  1: 0] nios_system_clock_2_out_byteenable;
  input            nios_system_clock_2_out_granted_sdram_0_s1;
  input            nios_system_clock_2_out_qualified_request_sdram_0_s1;
  input            nios_system_clock_2_out_read;
  input            nios_system_clock_2_out_read_data_valid_sdram_0_s1;
  input            nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register;
  input            nios_system_clock_2_out_requests_sdram_0_s1;
  input            nios_system_clock_2_out_write;
  input   [ 15: 0] nios_system_clock_2_out_writedata;
  input            reset_n;
  input   [ 15: 0] sdram_0_s1_readdata_from_sa;
  input            sdram_0_s1_waitrequest_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 22: 0] nios_system_clock_2_out_address_last_time;
  wire    [ 22: 0] nios_system_clock_2_out_address_to_slave;
  reg     [  1: 0] nios_system_clock_2_out_byteenable_last_time;
  reg              nios_system_clock_2_out_read_last_time;
  wire    [ 15: 0] nios_system_clock_2_out_readdata;
  wire             nios_system_clock_2_out_reset_n;
  wire             nios_system_clock_2_out_run;
  wire             nios_system_clock_2_out_waitrequest;
  reg              nios_system_clock_2_out_write_last_time;
  reg     [ 15: 0] nios_system_clock_2_out_writedata_last_time;
  wire             r_3;
  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (nios_system_clock_2_out_qualified_request_sdram_0_s1 | nios_system_clock_2_out_read_data_valid_sdram_0_s1 | ~nios_system_clock_2_out_requests_sdram_0_s1) & (nios_system_clock_2_out_granted_sdram_0_s1 | ~nios_system_clock_2_out_qualified_request_sdram_0_s1) & ((~nios_system_clock_2_out_qualified_request_sdram_0_s1 | ~nios_system_clock_2_out_read | (nios_system_clock_2_out_read_data_valid_sdram_0_s1 & nios_system_clock_2_out_read))) & ((~nios_system_clock_2_out_qualified_request_sdram_0_s1 | ~(nios_system_clock_2_out_read | nios_system_clock_2_out_write) | (1 & ~sdram_0_s1_waitrequest_from_sa & (nios_system_clock_2_out_read | nios_system_clock_2_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_2_out_run = r_3;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_2_out_address_to_slave = nios_system_clock_2_out_address;

  //nios_system_clock_2/out readdata mux, which is an e_mux
  assign nios_system_clock_2_out_readdata = sdram_0_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_2_out_waitrequest = ~nios_system_clock_2_out_run;

  //nios_system_clock_2_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_2_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_2_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_2_out_address_last_time <= 0;
      else 
        nios_system_clock_2_out_address_last_time <= nios_system_clock_2_out_address;
    end


  //nios_system_clock_2/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_2_out_waitrequest & (nios_system_clock_2_out_read | nios_system_clock_2_out_write);
    end


  //nios_system_clock_2_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_2_out_address != nios_system_clock_2_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_2_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_2_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_2_out_byteenable_last_time <= 0;
      else 
        nios_system_clock_2_out_byteenable_last_time <= nios_system_clock_2_out_byteenable;
    end


  //nios_system_clock_2_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_2_out_byteenable != nios_system_clock_2_out_byteenable_last_time))
        begin
          $write("%0d ns: nios_system_clock_2_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_2_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_2_out_read_last_time <= 0;
      else 
        nios_system_clock_2_out_read_last_time <= nios_system_clock_2_out_read;
    end


  //nios_system_clock_2_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_2_out_read != nios_system_clock_2_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_2_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_2_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_2_out_write_last_time <= 0;
      else 
        nios_system_clock_2_out_write_last_time <= nios_system_clock_2_out_write;
    end


  //nios_system_clock_2_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_2_out_write != nios_system_clock_2_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_2_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_2_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_2_out_writedata_last_time <= 0;
      else 
        nios_system_clock_2_out_writedata_last_time <= nios_system_clock_2_out_writedata;
    end


  //nios_system_clock_2_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_2_out_writedata != nios_system_clock_2_out_writedata_last_time) & nios_system_clock_2_out_write)
        begin
          $write("%0d ns: nios_system_clock_2_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_3_in_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_0_data_master_address_to_slave,
                                            cpu_0_data_master_byteenable,
                                            cpu_0_data_master_dbs_address,
                                            cpu_0_data_master_dbs_write_16,
                                            cpu_0_data_master_latency_counter,
                                            cpu_0_data_master_read,
                                            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                            cpu_0_data_master_write,
                                            nios_system_clock_3_in_endofpacket,
                                            nios_system_clock_3_in_readdata,
                                            nios_system_clock_3_in_waitrequest,
                                            reset_n,

                                           // outputs:
                                            cpu_0_data_master_byteenable_nios_system_clock_3_in,
                                            cpu_0_data_master_granted_nios_system_clock_3_in,
                                            cpu_0_data_master_qualified_request_nios_system_clock_3_in,
                                            cpu_0_data_master_read_data_valid_nios_system_clock_3_in,
                                            cpu_0_data_master_requests_nios_system_clock_3_in,
                                            d1_nios_system_clock_3_in_end_xfer,
                                            nios_system_clock_3_in_address,
                                            nios_system_clock_3_in_byteenable,
                                            nios_system_clock_3_in_endofpacket_from_sa,
                                            nios_system_clock_3_in_nativeaddress,
                                            nios_system_clock_3_in_read,
                                            nios_system_clock_3_in_readdata_from_sa,
                                            nios_system_clock_3_in_reset_n,
                                            nios_system_clock_3_in_waitrequest_from_sa,
                                            nios_system_clock_3_in_write,
                                            nios_system_clock_3_in_writedata
                                         )
;

  output  [  1: 0] cpu_0_data_master_byteenable_nios_system_clock_3_in;
  output           cpu_0_data_master_granted_nios_system_clock_3_in;
  output           cpu_0_data_master_qualified_request_nios_system_clock_3_in;
  output           cpu_0_data_master_read_data_valid_nios_system_clock_3_in;
  output           cpu_0_data_master_requests_nios_system_clock_3_in;
  output           d1_nios_system_clock_3_in_end_xfer;
  output  [ 22: 0] nios_system_clock_3_in_address;
  output  [  1: 0] nios_system_clock_3_in_byteenable;
  output           nios_system_clock_3_in_endofpacket_from_sa;
  output  [ 21: 0] nios_system_clock_3_in_nativeaddress;
  output           nios_system_clock_3_in_read;
  output  [ 15: 0] nios_system_clock_3_in_readdata_from_sa;
  output           nios_system_clock_3_in_reset_n;
  output           nios_system_clock_3_in_waitrequest_from_sa;
  output           nios_system_clock_3_in_write;
  output  [ 15: 0] nios_system_clock_3_in_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input   [  1: 0] cpu_0_data_master_dbs_address;
  input   [ 15: 0] cpu_0_data_master_dbs_write_16;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input            nios_system_clock_3_in_endofpacket;
  input   [ 15: 0] nios_system_clock_3_in_readdata;
  input            nios_system_clock_3_in_waitrequest;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire    [  1: 0] cpu_0_data_master_byteenable_nios_system_clock_3_in;
  wire    [  1: 0] cpu_0_data_master_byteenable_nios_system_clock_3_in_segment_0;
  wire    [  1: 0] cpu_0_data_master_byteenable_nios_system_clock_3_in_segment_1;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_nios_system_clock_3_in;
  wire             cpu_0_data_master_qualified_request_nios_system_clock_3_in;
  wire             cpu_0_data_master_read_data_valid_nios_system_clock_3_in;
  wire             cpu_0_data_master_requests_nios_system_clock_3_in;
  wire             cpu_0_data_master_saved_grant_nios_system_clock_3_in;
  reg              d1_nios_system_clock_3_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_3_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 22: 0] nios_system_clock_3_in_address;
  wire             nios_system_clock_3_in_allgrants;
  wire             nios_system_clock_3_in_allow_new_arb_cycle;
  wire             nios_system_clock_3_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_3_in_any_continuerequest;
  wire             nios_system_clock_3_in_arb_counter_enable;
  reg     [  2: 0] nios_system_clock_3_in_arb_share_counter;
  wire    [  2: 0] nios_system_clock_3_in_arb_share_counter_next_value;
  wire    [  2: 0] nios_system_clock_3_in_arb_share_set_values;
  wire             nios_system_clock_3_in_beginbursttransfer_internal;
  wire             nios_system_clock_3_in_begins_xfer;
  wire    [  1: 0] nios_system_clock_3_in_byteenable;
  wire             nios_system_clock_3_in_end_xfer;
  wire             nios_system_clock_3_in_endofpacket_from_sa;
  wire             nios_system_clock_3_in_firsttransfer;
  wire             nios_system_clock_3_in_grant_vector;
  wire             nios_system_clock_3_in_in_a_read_cycle;
  wire             nios_system_clock_3_in_in_a_write_cycle;
  wire             nios_system_clock_3_in_master_qreq_vector;
  wire    [ 21: 0] nios_system_clock_3_in_nativeaddress;
  wire             nios_system_clock_3_in_non_bursting_master_requests;
  wire             nios_system_clock_3_in_read;
  wire    [ 15: 0] nios_system_clock_3_in_readdata_from_sa;
  reg              nios_system_clock_3_in_reg_firsttransfer;
  wire             nios_system_clock_3_in_reset_n;
  reg              nios_system_clock_3_in_slavearbiterlockenable;
  wire             nios_system_clock_3_in_slavearbiterlockenable2;
  wire             nios_system_clock_3_in_unreg_firsttransfer;
  wire             nios_system_clock_3_in_waitrequest_from_sa;
  wire             nios_system_clock_3_in_waits_for_read;
  wire             nios_system_clock_3_in_waits_for_write;
  wire             nios_system_clock_3_in_write;
  wire    [ 15: 0] nios_system_clock_3_in_writedata;
  wire             wait_for_nios_system_clock_3_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_3_in_end_xfer;
    end


  assign nios_system_clock_3_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_nios_system_clock_3_in));
  //assign nios_system_clock_3_in_readdata_from_sa = nios_system_clock_3_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_3_in_readdata_from_sa = nios_system_clock_3_in_readdata;

  assign cpu_0_data_master_requests_nios_system_clock_3_in = ({cpu_0_data_master_address_to_slave[24 : 23] , 23'b0} == 25'h800000) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //assign nios_system_clock_3_in_waitrequest_from_sa = nios_system_clock_3_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_3_in_waitrequest_from_sa = nios_system_clock_3_in_waitrequest;

  //nios_system_clock_3_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_3_in_arb_share_set_values = (cpu_0_data_master_granted_nios_system_clock_3_in)? 2 :
    1;

  //nios_system_clock_3_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_3_in_non_bursting_master_requests = cpu_0_data_master_requests_nios_system_clock_3_in;

  //nios_system_clock_3_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_3_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_3_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_3_in_arb_share_counter_next_value = nios_system_clock_3_in_firsttransfer ? (nios_system_clock_3_in_arb_share_set_values - 1) : |nios_system_clock_3_in_arb_share_counter ? (nios_system_clock_3_in_arb_share_counter - 1) : 0;

  //nios_system_clock_3_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_3_in_allgrants = |nios_system_clock_3_in_grant_vector;

  //nios_system_clock_3_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_3_in_end_xfer = ~(nios_system_clock_3_in_waits_for_read | nios_system_clock_3_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_3_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_3_in = nios_system_clock_3_in_end_xfer & (~nios_system_clock_3_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_3_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_3_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_3_in & nios_system_clock_3_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_3_in & ~nios_system_clock_3_in_non_bursting_master_requests);

  //nios_system_clock_3_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_3_in_arb_share_counter <= 0;
      else if (nios_system_clock_3_in_arb_counter_enable)
          nios_system_clock_3_in_arb_share_counter <= nios_system_clock_3_in_arb_share_counter_next_value;
    end


  //nios_system_clock_3_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_3_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_3_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_3_in) | (end_xfer_arb_share_counter_term_nios_system_clock_3_in & ~nios_system_clock_3_in_non_bursting_master_requests))
          nios_system_clock_3_in_slavearbiterlockenable <= |nios_system_clock_3_in_arb_share_counter_next_value;
    end


  //cpu_0/data_master nios_system_clock_3/in arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = nios_system_clock_3_in_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //nios_system_clock_3_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_3_in_slavearbiterlockenable2 = |nios_system_clock_3_in_arb_share_counter_next_value;

  //cpu_0/data_master nios_system_clock_3/in arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = nios_system_clock_3_in_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //nios_system_clock_3_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_3_in_any_continuerequest = 1;

  //cpu_0_data_master_continuerequest continued request, which is an e_assign
  assign cpu_0_data_master_continuerequest = 1;

  assign cpu_0_data_master_qualified_request_nios_system_clock_3_in = cpu_0_data_master_requests_nios_system_clock_3_in & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | ((!cpu_0_data_master_byteenable_nios_system_clock_3_in) & cpu_0_data_master_write));
  //local readdatavalid cpu_0_data_master_read_data_valid_nios_system_clock_3_in, which is an e_mux
  assign cpu_0_data_master_read_data_valid_nios_system_clock_3_in = cpu_0_data_master_granted_nios_system_clock_3_in & cpu_0_data_master_read & ~nios_system_clock_3_in_waits_for_read;

  //nios_system_clock_3_in_writedata mux, which is an e_mux
  assign nios_system_clock_3_in_writedata = cpu_0_data_master_dbs_write_16;

  //assign nios_system_clock_3_in_endofpacket_from_sa = nios_system_clock_3_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_3_in_endofpacket_from_sa = nios_system_clock_3_in_endofpacket;

  //master is always granted when requested
  assign cpu_0_data_master_granted_nios_system_clock_3_in = cpu_0_data_master_qualified_request_nios_system_clock_3_in;

  //cpu_0/data_master saved-grant nios_system_clock_3/in, which is an e_assign
  assign cpu_0_data_master_saved_grant_nios_system_clock_3_in = cpu_0_data_master_requests_nios_system_clock_3_in;

  //allow new arb cycle for nios_system_clock_3/in, which is an e_assign
  assign nios_system_clock_3_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_3_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_3_in_master_qreq_vector = 1;

  //nios_system_clock_3_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_3_in_reset_n = reset_n;

  //nios_system_clock_3_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_3_in_firsttransfer = nios_system_clock_3_in_begins_xfer ? nios_system_clock_3_in_unreg_firsttransfer : nios_system_clock_3_in_reg_firsttransfer;

  //nios_system_clock_3_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_3_in_unreg_firsttransfer = ~(nios_system_clock_3_in_slavearbiterlockenable & nios_system_clock_3_in_any_continuerequest);

  //nios_system_clock_3_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_3_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_3_in_begins_xfer)
          nios_system_clock_3_in_reg_firsttransfer <= nios_system_clock_3_in_unreg_firsttransfer;
    end


  //nios_system_clock_3_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_3_in_beginbursttransfer_internal = nios_system_clock_3_in_begins_xfer;

  //nios_system_clock_3_in_read assignment, which is an e_mux
  assign nios_system_clock_3_in_read = cpu_0_data_master_granted_nios_system_clock_3_in & cpu_0_data_master_read;

  //nios_system_clock_3_in_write assignment, which is an e_mux
  assign nios_system_clock_3_in_write = cpu_0_data_master_granted_nios_system_clock_3_in & cpu_0_data_master_write;

  //nios_system_clock_3_in_address mux, which is an e_mux
  assign nios_system_clock_3_in_address = {cpu_0_data_master_address_to_slave >> 2,
    cpu_0_data_master_dbs_address[1],
    {1 {1'b0}}};

  //slaveid nios_system_clock_3_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_3_in_nativeaddress = cpu_0_data_master_address_to_slave >> 2;

  //d1_nios_system_clock_3_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_3_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_3_in_end_xfer <= nios_system_clock_3_in_end_xfer;
    end


  //nios_system_clock_3_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_3_in_waits_for_read = nios_system_clock_3_in_in_a_read_cycle & nios_system_clock_3_in_waitrequest_from_sa;

  //nios_system_clock_3_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_3_in_in_a_read_cycle = cpu_0_data_master_granted_nios_system_clock_3_in & cpu_0_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_3_in_in_a_read_cycle;

  //nios_system_clock_3_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_3_in_waits_for_write = nios_system_clock_3_in_in_a_write_cycle & nios_system_clock_3_in_waitrequest_from_sa;

  //nios_system_clock_3_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_3_in_in_a_write_cycle = cpu_0_data_master_granted_nios_system_clock_3_in & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_3_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_3_in_counter = 0;
  //nios_system_clock_3_in_byteenable byte enable port mux, which is an e_mux
  assign nios_system_clock_3_in_byteenable = (cpu_0_data_master_granted_nios_system_clock_3_in)? cpu_0_data_master_byteenable_nios_system_clock_3_in :
    -1;

  assign {cpu_0_data_master_byteenable_nios_system_clock_3_in_segment_1,
cpu_0_data_master_byteenable_nios_system_clock_3_in_segment_0} = cpu_0_data_master_byteenable;
  assign cpu_0_data_master_byteenable_nios_system_clock_3_in = ((cpu_0_data_master_dbs_address[1] == 0))? cpu_0_data_master_byteenable_nios_system_clock_3_in_segment_0 :
    cpu_0_data_master_byteenable_nios_system_clock_3_in_segment_1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_3/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_3_out_arbitrator (
                                            // inputs:
                                             clk,
                                             d1_sdram_0_s1_end_xfer,
                                             nios_system_clock_3_out_address,
                                             nios_system_clock_3_out_byteenable,
                                             nios_system_clock_3_out_granted_sdram_0_s1,
                                             nios_system_clock_3_out_qualified_request_sdram_0_s1,
                                             nios_system_clock_3_out_read,
                                             nios_system_clock_3_out_read_data_valid_sdram_0_s1,
                                             nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register,
                                             nios_system_clock_3_out_requests_sdram_0_s1,
                                             nios_system_clock_3_out_write,
                                             nios_system_clock_3_out_writedata,
                                             reset_n,
                                             sdram_0_s1_readdata_from_sa,
                                             sdram_0_s1_waitrequest_from_sa,

                                            // outputs:
                                             nios_system_clock_3_out_address_to_slave,
                                             nios_system_clock_3_out_readdata,
                                             nios_system_clock_3_out_reset_n,
                                             nios_system_clock_3_out_waitrequest
                                          )
;

  output  [ 22: 0] nios_system_clock_3_out_address_to_slave;
  output  [ 15: 0] nios_system_clock_3_out_readdata;
  output           nios_system_clock_3_out_reset_n;
  output           nios_system_clock_3_out_waitrequest;
  input            clk;
  input            d1_sdram_0_s1_end_xfer;
  input   [ 22: 0] nios_system_clock_3_out_address;
  input   [  1: 0] nios_system_clock_3_out_byteenable;
  input            nios_system_clock_3_out_granted_sdram_0_s1;
  input            nios_system_clock_3_out_qualified_request_sdram_0_s1;
  input            nios_system_clock_3_out_read;
  input            nios_system_clock_3_out_read_data_valid_sdram_0_s1;
  input            nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register;
  input            nios_system_clock_3_out_requests_sdram_0_s1;
  input            nios_system_clock_3_out_write;
  input   [ 15: 0] nios_system_clock_3_out_writedata;
  input            reset_n;
  input   [ 15: 0] sdram_0_s1_readdata_from_sa;
  input            sdram_0_s1_waitrequest_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 22: 0] nios_system_clock_3_out_address_last_time;
  wire    [ 22: 0] nios_system_clock_3_out_address_to_slave;
  reg     [  1: 0] nios_system_clock_3_out_byteenable_last_time;
  reg              nios_system_clock_3_out_read_last_time;
  wire    [ 15: 0] nios_system_clock_3_out_readdata;
  wire             nios_system_clock_3_out_reset_n;
  wire             nios_system_clock_3_out_run;
  wire             nios_system_clock_3_out_waitrequest;
  reg              nios_system_clock_3_out_write_last_time;
  reg     [ 15: 0] nios_system_clock_3_out_writedata_last_time;
  wire             r_3;
  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (nios_system_clock_3_out_qualified_request_sdram_0_s1 | nios_system_clock_3_out_read_data_valid_sdram_0_s1 | ~nios_system_clock_3_out_requests_sdram_0_s1) & (nios_system_clock_3_out_granted_sdram_0_s1 | ~nios_system_clock_3_out_qualified_request_sdram_0_s1) & ((~nios_system_clock_3_out_qualified_request_sdram_0_s1 | ~nios_system_clock_3_out_read | (nios_system_clock_3_out_read_data_valid_sdram_0_s1 & nios_system_clock_3_out_read))) & ((~nios_system_clock_3_out_qualified_request_sdram_0_s1 | ~(nios_system_clock_3_out_read | nios_system_clock_3_out_write) | (1 & ~sdram_0_s1_waitrequest_from_sa & (nios_system_clock_3_out_read | nios_system_clock_3_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_3_out_run = r_3;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_3_out_address_to_slave = nios_system_clock_3_out_address;

  //nios_system_clock_3/out readdata mux, which is an e_mux
  assign nios_system_clock_3_out_readdata = sdram_0_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_3_out_waitrequest = ~nios_system_clock_3_out_run;

  //nios_system_clock_3_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_3_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_3_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_3_out_address_last_time <= 0;
      else 
        nios_system_clock_3_out_address_last_time <= nios_system_clock_3_out_address;
    end


  //nios_system_clock_3/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_3_out_waitrequest & (nios_system_clock_3_out_read | nios_system_clock_3_out_write);
    end


  //nios_system_clock_3_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_3_out_address != nios_system_clock_3_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_3_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_3_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_3_out_byteenable_last_time <= 0;
      else 
        nios_system_clock_3_out_byteenable_last_time <= nios_system_clock_3_out_byteenable;
    end


  //nios_system_clock_3_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_3_out_byteenable != nios_system_clock_3_out_byteenable_last_time))
        begin
          $write("%0d ns: nios_system_clock_3_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_3_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_3_out_read_last_time <= 0;
      else 
        nios_system_clock_3_out_read_last_time <= nios_system_clock_3_out_read;
    end


  //nios_system_clock_3_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_3_out_read != nios_system_clock_3_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_3_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_3_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_3_out_write_last_time <= 0;
      else 
        nios_system_clock_3_out_write_last_time <= nios_system_clock_3_out_write;
    end


  //nios_system_clock_3_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_3_out_write != nios_system_clock_3_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_3_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_3_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_3_out_writedata_last_time <= 0;
      else 
        nios_system_clock_3_out_writedata_last_time <= nios_system_clock_3_out_writedata;
    end


  //nios_system_clock_3_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_3_out_writedata != nios_system_clock_3_out_writedata_last_time) & nios_system_clock_3_out_write)
        begin
          $write("%0d ns: nios_system_clock_3_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_4_in_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_2_instruction_master_address_to_slave,
                                            cpu_2_instruction_master_dbs_address,
                                            cpu_2_instruction_master_latency_counter,
                                            cpu_2_instruction_master_read,
                                            cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                            nios_system_clock_4_in_endofpacket,
                                            nios_system_clock_4_in_readdata,
                                            nios_system_clock_4_in_waitrequest,
                                            reset_n,

                                           // outputs:
                                            cpu_2_instruction_master_granted_nios_system_clock_4_in,
                                            cpu_2_instruction_master_qualified_request_nios_system_clock_4_in,
                                            cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in,
                                            cpu_2_instruction_master_requests_nios_system_clock_4_in,
                                            d1_nios_system_clock_4_in_end_xfer,
                                            nios_system_clock_4_in_address,
                                            nios_system_clock_4_in_byteenable,
                                            nios_system_clock_4_in_endofpacket_from_sa,
                                            nios_system_clock_4_in_nativeaddress,
                                            nios_system_clock_4_in_read,
                                            nios_system_clock_4_in_readdata_from_sa,
                                            nios_system_clock_4_in_reset_n,
                                            nios_system_clock_4_in_waitrequest_from_sa,
                                            nios_system_clock_4_in_write
                                         )
;

  output           cpu_2_instruction_master_granted_nios_system_clock_4_in;
  output           cpu_2_instruction_master_qualified_request_nios_system_clock_4_in;
  output           cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in;
  output           cpu_2_instruction_master_requests_nios_system_clock_4_in;
  output           d1_nios_system_clock_4_in_end_xfer;
  output  [ 22: 0] nios_system_clock_4_in_address;
  output  [  1: 0] nios_system_clock_4_in_byteenable;
  output           nios_system_clock_4_in_endofpacket_from_sa;
  output  [ 21: 0] nios_system_clock_4_in_nativeaddress;
  output           nios_system_clock_4_in_read;
  output  [ 15: 0] nios_system_clock_4_in_readdata_from_sa;
  output           nios_system_clock_4_in_reset_n;
  output           nios_system_clock_4_in_waitrequest_from_sa;
  output           nios_system_clock_4_in_write;
  input            clk;
  input   [ 24: 0] cpu_2_instruction_master_address_to_slave;
  input   [  1: 0] cpu_2_instruction_master_dbs_address;
  input            cpu_2_instruction_master_latency_counter;
  input            cpu_2_instruction_master_read;
  input            cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            nios_system_clock_4_in_endofpacket;
  input   [ 15: 0] nios_system_clock_4_in_readdata;
  input            nios_system_clock_4_in_waitrequest;
  input            reset_n;

  wire             cpu_2_instruction_master_arbiterlock;
  wire             cpu_2_instruction_master_arbiterlock2;
  wire             cpu_2_instruction_master_continuerequest;
  wire             cpu_2_instruction_master_granted_nios_system_clock_4_in;
  wire             cpu_2_instruction_master_qualified_request_nios_system_clock_4_in;
  wire             cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in;
  wire             cpu_2_instruction_master_requests_nios_system_clock_4_in;
  wire             cpu_2_instruction_master_saved_grant_nios_system_clock_4_in;
  reg              d1_nios_system_clock_4_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_4_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 22: 0] nios_system_clock_4_in_address;
  wire             nios_system_clock_4_in_allgrants;
  wire             nios_system_clock_4_in_allow_new_arb_cycle;
  wire             nios_system_clock_4_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_4_in_any_continuerequest;
  wire             nios_system_clock_4_in_arb_counter_enable;
  reg     [  1: 0] nios_system_clock_4_in_arb_share_counter;
  wire    [  1: 0] nios_system_clock_4_in_arb_share_counter_next_value;
  wire    [  1: 0] nios_system_clock_4_in_arb_share_set_values;
  wire             nios_system_clock_4_in_beginbursttransfer_internal;
  wire             nios_system_clock_4_in_begins_xfer;
  wire    [  1: 0] nios_system_clock_4_in_byteenable;
  wire             nios_system_clock_4_in_end_xfer;
  wire             nios_system_clock_4_in_endofpacket_from_sa;
  wire             nios_system_clock_4_in_firsttransfer;
  wire             nios_system_clock_4_in_grant_vector;
  wire             nios_system_clock_4_in_in_a_read_cycle;
  wire             nios_system_clock_4_in_in_a_write_cycle;
  wire             nios_system_clock_4_in_master_qreq_vector;
  wire    [ 21: 0] nios_system_clock_4_in_nativeaddress;
  wire             nios_system_clock_4_in_non_bursting_master_requests;
  wire             nios_system_clock_4_in_read;
  wire    [ 15: 0] nios_system_clock_4_in_readdata_from_sa;
  reg              nios_system_clock_4_in_reg_firsttransfer;
  wire             nios_system_clock_4_in_reset_n;
  reg              nios_system_clock_4_in_slavearbiterlockenable;
  wire             nios_system_clock_4_in_slavearbiterlockenable2;
  wire             nios_system_clock_4_in_unreg_firsttransfer;
  wire             nios_system_clock_4_in_waitrequest_from_sa;
  wire             nios_system_clock_4_in_waits_for_read;
  wire             nios_system_clock_4_in_waits_for_write;
  wire             nios_system_clock_4_in_write;
  wire             wait_for_nios_system_clock_4_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_4_in_end_xfer;
    end


  assign nios_system_clock_4_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_2_instruction_master_qualified_request_nios_system_clock_4_in));
  //assign nios_system_clock_4_in_readdata_from_sa = nios_system_clock_4_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_4_in_readdata_from_sa = nios_system_clock_4_in_readdata;

  assign cpu_2_instruction_master_requests_nios_system_clock_4_in = (({cpu_2_instruction_master_address_to_slave[24 : 23] , 23'b0} == 25'h800000) & (cpu_2_instruction_master_read)) & cpu_2_instruction_master_read;
  //assign nios_system_clock_4_in_waitrequest_from_sa = nios_system_clock_4_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_4_in_waitrequest_from_sa = nios_system_clock_4_in_waitrequest;

  //nios_system_clock_4_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_4_in_arb_share_set_values = (cpu_2_instruction_master_granted_nios_system_clock_4_in)? 2 :
    1;

  //nios_system_clock_4_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_4_in_non_bursting_master_requests = cpu_2_instruction_master_requests_nios_system_clock_4_in;

  //nios_system_clock_4_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_4_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_4_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_4_in_arb_share_counter_next_value = nios_system_clock_4_in_firsttransfer ? (nios_system_clock_4_in_arb_share_set_values - 1) : |nios_system_clock_4_in_arb_share_counter ? (nios_system_clock_4_in_arb_share_counter - 1) : 0;

  //nios_system_clock_4_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_4_in_allgrants = |nios_system_clock_4_in_grant_vector;

  //nios_system_clock_4_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_4_in_end_xfer = ~(nios_system_clock_4_in_waits_for_read | nios_system_clock_4_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_4_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_4_in = nios_system_clock_4_in_end_xfer & (~nios_system_clock_4_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_4_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_4_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_4_in & nios_system_clock_4_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_4_in & ~nios_system_clock_4_in_non_bursting_master_requests);

  //nios_system_clock_4_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_4_in_arb_share_counter <= 0;
      else if (nios_system_clock_4_in_arb_counter_enable)
          nios_system_clock_4_in_arb_share_counter <= nios_system_clock_4_in_arb_share_counter_next_value;
    end


  //nios_system_clock_4_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_4_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_4_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_4_in) | (end_xfer_arb_share_counter_term_nios_system_clock_4_in & ~nios_system_clock_4_in_non_bursting_master_requests))
          nios_system_clock_4_in_slavearbiterlockenable <= |nios_system_clock_4_in_arb_share_counter_next_value;
    end


  //cpu_2/instruction_master nios_system_clock_4/in arbiterlock, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock = nios_system_clock_4_in_slavearbiterlockenable & cpu_2_instruction_master_continuerequest;

  //nios_system_clock_4_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_4_in_slavearbiterlockenable2 = |nios_system_clock_4_in_arb_share_counter_next_value;

  //cpu_2/instruction_master nios_system_clock_4/in arbiterlock2, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock2 = nios_system_clock_4_in_slavearbiterlockenable2 & cpu_2_instruction_master_continuerequest;

  //nios_system_clock_4_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_4_in_any_continuerequest = 1;

  //cpu_2_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_2_instruction_master_continuerequest = 1;

  assign cpu_2_instruction_master_qualified_request_nios_system_clock_4_in = cpu_2_instruction_master_requests_nios_system_clock_4_in & ~((cpu_2_instruction_master_read & ((cpu_2_instruction_master_latency_counter != 0) | (|cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))));
  //local readdatavalid cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in, which is an e_mux
  assign cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in = cpu_2_instruction_master_granted_nios_system_clock_4_in & cpu_2_instruction_master_read & ~nios_system_clock_4_in_waits_for_read;

  //assign nios_system_clock_4_in_endofpacket_from_sa = nios_system_clock_4_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_4_in_endofpacket_from_sa = nios_system_clock_4_in_endofpacket;

  //master is always granted when requested
  assign cpu_2_instruction_master_granted_nios_system_clock_4_in = cpu_2_instruction_master_qualified_request_nios_system_clock_4_in;

  //cpu_2/instruction_master saved-grant nios_system_clock_4/in, which is an e_assign
  assign cpu_2_instruction_master_saved_grant_nios_system_clock_4_in = cpu_2_instruction_master_requests_nios_system_clock_4_in;

  //allow new arb cycle for nios_system_clock_4/in, which is an e_assign
  assign nios_system_clock_4_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_4_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_4_in_master_qreq_vector = 1;

  //nios_system_clock_4_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_4_in_reset_n = reset_n;

  //nios_system_clock_4_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_4_in_firsttransfer = nios_system_clock_4_in_begins_xfer ? nios_system_clock_4_in_unreg_firsttransfer : nios_system_clock_4_in_reg_firsttransfer;

  //nios_system_clock_4_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_4_in_unreg_firsttransfer = ~(nios_system_clock_4_in_slavearbiterlockenable & nios_system_clock_4_in_any_continuerequest);

  //nios_system_clock_4_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_4_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_4_in_begins_xfer)
          nios_system_clock_4_in_reg_firsttransfer <= nios_system_clock_4_in_unreg_firsttransfer;
    end


  //nios_system_clock_4_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_4_in_beginbursttransfer_internal = nios_system_clock_4_in_begins_xfer;

  //nios_system_clock_4_in_read assignment, which is an e_mux
  assign nios_system_clock_4_in_read = cpu_2_instruction_master_granted_nios_system_clock_4_in & cpu_2_instruction_master_read;

  //nios_system_clock_4_in_write assignment, which is an e_mux
  assign nios_system_clock_4_in_write = 0;

  //nios_system_clock_4_in_address mux, which is an e_mux
  assign nios_system_clock_4_in_address = {cpu_2_instruction_master_address_to_slave >> 2,
    cpu_2_instruction_master_dbs_address[1],
    {1 {1'b0}}};

  //slaveid nios_system_clock_4_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_4_in_nativeaddress = cpu_2_instruction_master_address_to_slave >> 2;

  //d1_nios_system_clock_4_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_4_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_4_in_end_xfer <= nios_system_clock_4_in_end_xfer;
    end


  //nios_system_clock_4_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_4_in_waits_for_read = nios_system_clock_4_in_in_a_read_cycle & nios_system_clock_4_in_waitrequest_from_sa;

  //nios_system_clock_4_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_4_in_in_a_read_cycle = cpu_2_instruction_master_granted_nios_system_clock_4_in & cpu_2_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_4_in_in_a_read_cycle;

  //nios_system_clock_4_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_4_in_waits_for_write = nios_system_clock_4_in_in_a_write_cycle & nios_system_clock_4_in_waitrequest_from_sa;

  //nios_system_clock_4_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_4_in_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_4_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_4_in_counter = 0;
  //nios_system_clock_4_in_byteenable byte enable port mux, which is an e_mux
  assign nios_system_clock_4_in_byteenable = -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_4/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_4_out_arbitrator (
                                            // inputs:
                                             clk,
                                             d1_sdram_0_s1_end_xfer,
                                             nios_system_clock_4_out_address,
                                             nios_system_clock_4_out_byteenable,
                                             nios_system_clock_4_out_granted_sdram_0_s1,
                                             nios_system_clock_4_out_qualified_request_sdram_0_s1,
                                             nios_system_clock_4_out_read,
                                             nios_system_clock_4_out_read_data_valid_sdram_0_s1,
                                             nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register,
                                             nios_system_clock_4_out_requests_sdram_0_s1,
                                             nios_system_clock_4_out_write,
                                             nios_system_clock_4_out_writedata,
                                             reset_n,
                                             sdram_0_s1_readdata_from_sa,
                                             sdram_0_s1_waitrequest_from_sa,

                                            // outputs:
                                             nios_system_clock_4_out_address_to_slave,
                                             nios_system_clock_4_out_readdata,
                                             nios_system_clock_4_out_reset_n,
                                             nios_system_clock_4_out_waitrequest
                                          )
;

  output  [ 22: 0] nios_system_clock_4_out_address_to_slave;
  output  [ 15: 0] nios_system_clock_4_out_readdata;
  output           nios_system_clock_4_out_reset_n;
  output           nios_system_clock_4_out_waitrequest;
  input            clk;
  input            d1_sdram_0_s1_end_xfer;
  input   [ 22: 0] nios_system_clock_4_out_address;
  input   [  1: 0] nios_system_clock_4_out_byteenable;
  input            nios_system_clock_4_out_granted_sdram_0_s1;
  input            nios_system_clock_4_out_qualified_request_sdram_0_s1;
  input            nios_system_clock_4_out_read;
  input            nios_system_clock_4_out_read_data_valid_sdram_0_s1;
  input            nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register;
  input            nios_system_clock_4_out_requests_sdram_0_s1;
  input            nios_system_clock_4_out_write;
  input   [ 15: 0] nios_system_clock_4_out_writedata;
  input            reset_n;
  input   [ 15: 0] sdram_0_s1_readdata_from_sa;
  input            sdram_0_s1_waitrequest_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 22: 0] nios_system_clock_4_out_address_last_time;
  wire    [ 22: 0] nios_system_clock_4_out_address_to_slave;
  reg     [  1: 0] nios_system_clock_4_out_byteenable_last_time;
  reg              nios_system_clock_4_out_read_last_time;
  wire    [ 15: 0] nios_system_clock_4_out_readdata;
  wire             nios_system_clock_4_out_reset_n;
  wire             nios_system_clock_4_out_run;
  wire             nios_system_clock_4_out_waitrequest;
  reg              nios_system_clock_4_out_write_last_time;
  reg     [ 15: 0] nios_system_clock_4_out_writedata_last_time;
  wire             r_3;
  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (nios_system_clock_4_out_qualified_request_sdram_0_s1 | nios_system_clock_4_out_read_data_valid_sdram_0_s1 | ~nios_system_clock_4_out_requests_sdram_0_s1) & (nios_system_clock_4_out_granted_sdram_0_s1 | ~nios_system_clock_4_out_qualified_request_sdram_0_s1) & ((~nios_system_clock_4_out_qualified_request_sdram_0_s1 | ~nios_system_clock_4_out_read | (nios_system_clock_4_out_read_data_valid_sdram_0_s1 & nios_system_clock_4_out_read))) & ((~nios_system_clock_4_out_qualified_request_sdram_0_s1 | ~(nios_system_clock_4_out_read | nios_system_clock_4_out_write) | (1 & ~sdram_0_s1_waitrequest_from_sa & (nios_system_clock_4_out_read | nios_system_clock_4_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_4_out_run = r_3;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_4_out_address_to_slave = nios_system_clock_4_out_address;

  //nios_system_clock_4/out readdata mux, which is an e_mux
  assign nios_system_clock_4_out_readdata = sdram_0_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_4_out_waitrequest = ~nios_system_clock_4_out_run;

  //nios_system_clock_4_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_4_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_4_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_4_out_address_last_time <= 0;
      else 
        nios_system_clock_4_out_address_last_time <= nios_system_clock_4_out_address;
    end


  //nios_system_clock_4/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_4_out_waitrequest & (nios_system_clock_4_out_read | nios_system_clock_4_out_write);
    end


  //nios_system_clock_4_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_4_out_address != nios_system_clock_4_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_4_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_4_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_4_out_byteenable_last_time <= 0;
      else 
        nios_system_clock_4_out_byteenable_last_time <= nios_system_clock_4_out_byteenable;
    end


  //nios_system_clock_4_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_4_out_byteenable != nios_system_clock_4_out_byteenable_last_time))
        begin
          $write("%0d ns: nios_system_clock_4_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_4_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_4_out_read_last_time <= 0;
      else 
        nios_system_clock_4_out_read_last_time <= nios_system_clock_4_out_read;
    end


  //nios_system_clock_4_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_4_out_read != nios_system_clock_4_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_4_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_4_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_4_out_write_last_time <= 0;
      else 
        nios_system_clock_4_out_write_last_time <= nios_system_clock_4_out_write;
    end


  //nios_system_clock_4_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_4_out_write != nios_system_clock_4_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_4_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_4_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_4_out_writedata_last_time <= 0;
      else 
        nios_system_clock_4_out_writedata_last_time <= nios_system_clock_4_out_writedata;
    end


  //nios_system_clock_4_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_4_out_writedata != nios_system_clock_4_out_writedata_last_time) & nios_system_clock_4_out_write)
        begin
          $write("%0d ns: nios_system_clock_4_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_5_in_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_2_data_master_address_to_slave,
                                            cpu_2_data_master_byteenable,
                                            cpu_2_data_master_dbs_address,
                                            cpu_2_data_master_dbs_write_16,
                                            cpu_2_data_master_latency_counter,
                                            cpu_2_data_master_read,
                                            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                            cpu_2_data_master_write,
                                            nios_system_clock_5_in_endofpacket,
                                            nios_system_clock_5_in_readdata,
                                            nios_system_clock_5_in_waitrequest,
                                            reset_n,

                                           // outputs:
                                            cpu_2_data_master_byteenable_nios_system_clock_5_in,
                                            cpu_2_data_master_granted_nios_system_clock_5_in,
                                            cpu_2_data_master_qualified_request_nios_system_clock_5_in,
                                            cpu_2_data_master_read_data_valid_nios_system_clock_5_in,
                                            cpu_2_data_master_requests_nios_system_clock_5_in,
                                            d1_nios_system_clock_5_in_end_xfer,
                                            nios_system_clock_5_in_address,
                                            nios_system_clock_5_in_byteenable,
                                            nios_system_clock_5_in_endofpacket_from_sa,
                                            nios_system_clock_5_in_nativeaddress,
                                            nios_system_clock_5_in_read,
                                            nios_system_clock_5_in_readdata_from_sa,
                                            nios_system_clock_5_in_reset_n,
                                            nios_system_clock_5_in_waitrequest_from_sa,
                                            nios_system_clock_5_in_write,
                                            nios_system_clock_5_in_writedata
                                         )
;

  output  [  1: 0] cpu_2_data_master_byteenable_nios_system_clock_5_in;
  output           cpu_2_data_master_granted_nios_system_clock_5_in;
  output           cpu_2_data_master_qualified_request_nios_system_clock_5_in;
  output           cpu_2_data_master_read_data_valid_nios_system_clock_5_in;
  output           cpu_2_data_master_requests_nios_system_clock_5_in;
  output           d1_nios_system_clock_5_in_end_xfer;
  output  [ 22: 0] nios_system_clock_5_in_address;
  output  [  1: 0] nios_system_clock_5_in_byteenable;
  output           nios_system_clock_5_in_endofpacket_from_sa;
  output  [ 21: 0] nios_system_clock_5_in_nativeaddress;
  output           nios_system_clock_5_in_read;
  output  [ 15: 0] nios_system_clock_5_in_readdata_from_sa;
  output           nios_system_clock_5_in_reset_n;
  output           nios_system_clock_5_in_waitrequest_from_sa;
  output           nios_system_clock_5_in_write;
  output  [ 15: 0] nios_system_clock_5_in_writedata;
  input            clk;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input   [  3: 0] cpu_2_data_master_byteenable;
  input   [  1: 0] cpu_2_data_master_dbs_address;
  input   [ 15: 0] cpu_2_data_master_dbs_write_16;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input            nios_system_clock_5_in_endofpacket;
  input   [ 15: 0] nios_system_clock_5_in_readdata;
  input            nios_system_clock_5_in_waitrequest;
  input            reset_n;

  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire    [  1: 0] cpu_2_data_master_byteenable_nios_system_clock_5_in;
  wire    [  1: 0] cpu_2_data_master_byteenable_nios_system_clock_5_in_segment_0;
  wire    [  1: 0] cpu_2_data_master_byteenable_nios_system_clock_5_in_segment_1;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_nios_system_clock_5_in;
  wire             cpu_2_data_master_qualified_request_nios_system_clock_5_in;
  wire             cpu_2_data_master_read_data_valid_nios_system_clock_5_in;
  wire             cpu_2_data_master_requests_nios_system_clock_5_in;
  wire             cpu_2_data_master_saved_grant_nios_system_clock_5_in;
  reg              d1_nios_system_clock_5_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_5_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 22: 0] nios_system_clock_5_in_address;
  wire             nios_system_clock_5_in_allgrants;
  wire             nios_system_clock_5_in_allow_new_arb_cycle;
  wire             nios_system_clock_5_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_5_in_any_continuerequest;
  wire             nios_system_clock_5_in_arb_counter_enable;
  reg     [  2: 0] nios_system_clock_5_in_arb_share_counter;
  wire    [  2: 0] nios_system_clock_5_in_arb_share_counter_next_value;
  wire    [  2: 0] nios_system_clock_5_in_arb_share_set_values;
  wire             nios_system_clock_5_in_beginbursttransfer_internal;
  wire             nios_system_clock_5_in_begins_xfer;
  wire    [  1: 0] nios_system_clock_5_in_byteenable;
  wire             nios_system_clock_5_in_end_xfer;
  wire             nios_system_clock_5_in_endofpacket_from_sa;
  wire             nios_system_clock_5_in_firsttransfer;
  wire             nios_system_clock_5_in_grant_vector;
  wire             nios_system_clock_5_in_in_a_read_cycle;
  wire             nios_system_clock_5_in_in_a_write_cycle;
  wire             nios_system_clock_5_in_master_qreq_vector;
  wire    [ 21: 0] nios_system_clock_5_in_nativeaddress;
  wire             nios_system_clock_5_in_non_bursting_master_requests;
  wire             nios_system_clock_5_in_read;
  wire    [ 15: 0] nios_system_clock_5_in_readdata_from_sa;
  reg              nios_system_clock_5_in_reg_firsttransfer;
  wire             nios_system_clock_5_in_reset_n;
  reg              nios_system_clock_5_in_slavearbiterlockenable;
  wire             nios_system_clock_5_in_slavearbiterlockenable2;
  wire             nios_system_clock_5_in_unreg_firsttransfer;
  wire             nios_system_clock_5_in_waitrequest_from_sa;
  wire             nios_system_clock_5_in_waits_for_read;
  wire             nios_system_clock_5_in_waits_for_write;
  wire             nios_system_clock_5_in_write;
  wire    [ 15: 0] nios_system_clock_5_in_writedata;
  wire             wait_for_nios_system_clock_5_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_5_in_end_xfer;
    end


  assign nios_system_clock_5_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_2_data_master_qualified_request_nios_system_clock_5_in));
  //assign nios_system_clock_5_in_readdata_from_sa = nios_system_clock_5_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_5_in_readdata_from_sa = nios_system_clock_5_in_readdata;

  assign cpu_2_data_master_requests_nios_system_clock_5_in = ({cpu_2_data_master_address_to_slave[24 : 23] , 23'b0} == 25'h800000) & (cpu_2_data_master_read | cpu_2_data_master_write);
  //assign nios_system_clock_5_in_waitrequest_from_sa = nios_system_clock_5_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_5_in_waitrequest_from_sa = nios_system_clock_5_in_waitrequest;

  //nios_system_clock_5_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_5_in_arb_share_set_values = (cpu_2_data_master_granted_nios_system_clock_5_in)? 2 :
    1;

  //nios_system_clock_5_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_5_in_non_bursting_master_requests = cpu_2_data_master_requests_nios_system_clock_5_in;

  //nios_system_clock_5_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_5_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_5_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_5_in_arb_share_counter_next_value = nios_system_clock_5_in_firsttransfer ? (nios_system_clock_5_in_arb_share_set_values - 1) : |nios_system_clock_5_in_arb_share_counter ? (nios_system_clock_5_in_arb_share_counter - 1) : 0;

  //nios_system_clock_5_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_5_in_allgrants = |nios_system_clock_5_in_grant_vector;

  //nios_system_clock_5_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_5_in_end_xfer = ~(nios_system_clock_5_in_waits_for_read | nios_system_clock_5_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_5_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_5_in = nios_system_clock_5_in_end_xfer & (~nios_system_clock_5_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_5_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_5_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_5_in & nios_system_clock_5_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_5_in & ~nios_system_clock_5_in_non_bursting_master_requests);

  //nios_system_clock_5_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_5_in_arb_share_counter <= 0;
      else if (nios_system_clock_5_in_arb_counter_enable)
          nios_system_clock_5_in_arb_share_counter <= nios_system_clock_5_in_arb_share_counter_next_value;
    end


  //nios_system_clock_5_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_5_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_5_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_5_in) | (end_xfer_arb_share_counter_term_nios_system_clock_5_in & ~nios_system_clock_5_in_non_bursting_master_requests))
          nios_system_clock_5_in_slavearbiterlockenable <= |nios_system_clock_5_in_arb_share_counter_next_value;
    end


  //cpu_2/data_master nios_system_clock_5/in arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = nios_system_clock_5_in_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //nios_system_clock_5_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_5_in_slavearbiterlockenable2 = |nios_system_clock_5_in_arb_share_counter_next_value;

  //cpu_2/data_master nios_system_clock_5/in arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = nios_system_clock_5_in_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //nios_system_clock_5_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_5_in_any_continuerequest = 1;

  //cpu_2_data_master_continuerequest continued request, which is an e_assign
  assign cpu_2_data_master_continuerequest = 1;

  assign cpu_2_data_master_qualified_request_nios_system_clock_5_in = cpu_2_data_master_requests_nios_system_clock_5_in & ~((cpu_2_data_master_read & ((cpu_2_data_master_latency_counter != 0) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | ((!cpu_2_data_master_byteenable_nios_system_clock_5_in) & cpu_2_data_master_write));
  //local readdatavalid cpu_2_data_master_read_data_valid_nios_system_clock_5_in, which is an e_mux
  assign cpu_2_data_master_read_data_valid_nios_system_clock_5_in = cpu_2_data_master_granted_nios_system_clock_5_in & cpu_2_data_master_read & ~nios_system_clock_5_in_waits_for_read;

  //nios_system_clock_5_in_writedata mux, which is an e_mux
  assign nios_system_clock_5_in_writedata = cpu_2_data_master_dbs_write_16;

  //assign nios_system_clock_5_in_endofpacket_from_sa = nios_system_clock_5_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_5_in_endofpacket_from_sa = nios_system_clock_5_in_endofpacket;

  //master is always granted when requested
  assign cpu_2_data_master_granted_nios_system_clock_5_in = cpu_2_data_master_qualified_request_nios_system_clock_5_in;

  //cpu_2/data_master saved-grant nios_system_clock_5/in, which is an e_assign
  assign cpu_2_data_master_saved_grant_nios_system_clock_5_in = cpu_2_data_master_requests_nios_system_clock_5_in;

  //allow new arb cycle for nios_system_clock_5/in, which is an e_assign
  assign nios_system_clock_5_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_5_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_5_in_master_qreq_vector = 1;

  //nios_system_clock_5_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_5_in_reset_n = reset_n;

  //nios_system_clock_5_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_5_in_firsttransfer = nios_system_clock_5_in_begins_xfer ? nios_system_clock_5_in_unreg_firsttransfer : nios_system_clock_5_in_reg_firsttransfer;

  //nios_system_clock_5_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_5_in_unreg_firsttransfer = ~(nios_system_clock_5_in_slavearbiterlockenable & nios_system_clock_5_in_any_continuerequest);

  //nios_system_clock_5_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_5_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_5_in_begins_xfer)
          nios_system_clock_5_in_reg_firsttransfer <= nios_system_clock_5_in_unreg_firsttransfer;
    end


  //nios_system_clock_5_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_5_in_beginbursttransfer_internal = nios_system_clock_5_in_begins_xfer;

  //nios_system_clock_5_in_read assignment, which is an e_mux
  assign nios_system_clock_5_in_read = cpu_2_data_master_granted_nios_system_clock_5_in & cpu_2_data_master_read;

  //nios_system_clock_5_in_write assignment, which is an e_mux
  assign nios_system_clock_5_in_write = cpu_2_data_master_granted_nios_system_clock_5_in & cpu_2_data_master_write;

  //nios_system_clock_5_in_address mux, which is an e_mux
  assign nios_system_clock_5_in_address = {cpu_2_data_master_address_to_slave >> 2,
    cpu_2_data_master_dbs_address[1],
    {1 {1'b0}}};

  //slaveid nios_system_clock_5_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_5_in_nativeaddress = cpu_2_data_master_address_to_slave >> 2;

  //d1_nios_system_clock_5_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_5_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_5_in_end_xfer <= nios_system_clock_5_in_end_xfer;
    end


  //nios_system_clock_5_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_5_in_waits_for_read = nios_system_clock_5_in_in_a_read_cycle & nios_system_clock_5_in_waitrequest_from_sa;

  //nios_system_clock_5_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_5_in_in_a_read_cycle = cpu_2_data_master_granted_nios_system_clock_5_in & cpu_2_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_5_in_in_a_read_cycle;

  //nios_system_clock_5_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_5_in_waits_for_write = nios_system_clock_5_in_in_a_write_cycle & nios_system_clock_5_in_waitrequest_from_sa;

  //nios_system_clock_5_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_5_in_in_a_write_cycle = cpu_2_data_master_granted_nios_system_clock_5_in & cpu_2_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_5_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_5_in_counter = 0;
  //nios_system_clock_5_in_byteenable byte enable port mux, which is an e_mux
  assign nios_system_clock_5_in_byteenable = (cpu_2_data_master_granted_nios_system_clock_5_in)? cpu_2_data_master_byteenable_nios_system_clock_5_in :
    -1;

  assign {cpu_2_data_master_byteenable_nios_system_clock_5_in_segment_1,
cpu_2_data_master_byteenable_nios_system_clock_5_in_segment_0} = cpu_2_data_master_byteenable;
  assign cpu_2_data_master_byteenable_nios_system_clock_5_in = ((cpu_2_data_master_dbs_address[1] == 0))? cpu_2_data_master_byteenable_nios_system_clock_5_in_segment_0 :
    cpu_2_data_master_byteenable_nios_system_clock_5_in_segment_1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_5/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_5_out_arbitrator (
                                            // inputs:
                                             clk,
                                             d1_sdram_0_s1_end_xfer,
                                             nios_system_clock_5_out_address,
                                             nios_system_clock_5_out_byteenable,
                                             nios_system_clock_5_out_granted_sdram_0_s1,
                                             nios_system_clock_5_out_qualified_request_sdram_0_s1,
                                             nios_system_clock_5_out_read,
                                             nios_system_clock_5_out_read_data_valid_sdram_0_s1,
                                             nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register,
                                             nios_system_clock_5_out_requests_sdram_0_s1,
                                             nios_system_clock_5_out_write,
                                             nios_system_clock_5_out_writedata,
                                             reset_n,
                                             sdram_0_s1_readdata_from_sa,
                                             sdram_0_s1_waitrequest_from_sa,

                                            // outputs:
                                             nios_system_clock_5_out_address_to_slave,
                                             nios_system_clock_5_out_readdata,
                                             nios_system_clock_5_out_reset_n,
                                             nios_system_clock_5_out_waitrequest
                                          )
;

  output  [ 22: 0] nios_system_clock_5_out_address_to_slave;
  output  [ 15: 0] nios_system_clock_5_out_readdata;
  output           nios_system_clock_5_out_reset_n;
  output           nios_system_clock_5_out_waitrequest;
  input            clk;
  input            d1_sdram_0_s1_end_xfer;
  input   [ 22: 0] nios_system_clock_5_out_address;
  input   [  1: 0] nios_system_clock_5_out_byteenable;
  input            nios_system_clock_5_out_granted_sdram_0_s1;
  input            nios_system_clock_5_out_qualified_request_sdram_0_s1;
  input            nios_system_clock_5_out_read;
  input            nios_system_clock_5_out_read_data_valid_sdram_0_s1;
  input            nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register;
  input            nios_system_clock_5_out_requests_sdram_0_s1;
  input            nios_system_clock_5_out_write;
  input   [ 15: 0] nios_system_clock_5_out_writedata;
  input            reset_n;
  input   [ 15: 0] sdram_0_s1_readdata_from_sa;
  input            sdram_0_s1_waitrequest_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 22: 0] nios_system_clock_5_out_address_last_time;
  wire    [ 22: 0] nios_system_clock_5_out_address_to_slave;
  reg     [  1: 0] nios_system_clock_5_out_byteenable_last_time;
  reg              nios_system_clock_5_out_read_last_time;
  wire    [ 15: 0] nios_system_clock_5_out_readdata;
  wire             nios_system_clock_5_out_reset_n;
  wire             nios_system_clock_5_out_run;
  wire             nios_system_clock_5_out_waitrequest;
  reg              nios_system_clock_5_out_write_last_time;
  reg     [ 15: 0] nios_system_clock_5_out_writedata_last_time;
  wire             r_3;
  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (nios_system_clock_5_out_qualified_request_sdram_0_s1 | nios_system_clock_5_out_read_data_valid_sdram_0_s1 | ~nios_system_clock_5_out_requests_sdram_0_s1) & (nios_system_clock_5_out_granted_sdram_0_s1 | ~nios_system_clock_5_out_qualified_request_sdram_0_s1) & ((~nios_system_clock_5_out_qualified_request_sdram_0_s1 | ~nios_system_clock_5_out_read | (nios_system_clock_5_out_read_data_valid_sdram_0_s1 & nios_system_clock_5_out_read))) & ((~nios_system_clock_5_out_qualified_request_sdram_0_s1 | ~(nios_system_clock_5_out_read | nios_system_clock_5_out_write) | (1 & ~sdram_0_s1_waitrequest_from_sa & (nios_system_clock_5_out_read | nios_system_clock_5_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_5_out_run = r_3;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_5_out_address_to_slave = nios_system_clock_5_out_address;

  //nios_system_clock_5/out readdata mux, which is an e_mux
  assign nios_system_clock_5_out_readdata = sdram_0_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_5_out_waitrequest = ~nios_system_clock_5_out_run;

  //nios_system_clock_5_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_5_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_5_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_5_out_address_last_time <= 0;
      else 
        nios_system_clock_5_out_address_last_time <= nios_system_clock_5_out_address;
    end


  //nios_system_clock_5/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_5_out_waitrequest & (nios_system_clock_5_out_read | nios_system_clock_5_out_write);
    end


  //nios_system_clock_5_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_5_out_address != nios_system_clock_5_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_5_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_5_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_5_out_byteenable_last_time <= 0;
      else 
        nios_system_clock_5_out_byteenable_last_time <= nios_system_clock_5_out_byteenable;
    end


  //nios_system_clock_5_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_5_out_byteenable != nios_system_clock_5_out_byteenable_last_time))
        begin
          $write("%0d ns: nios_system_clock_5_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_5_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_5_out_read_last_time <= 0;
      else 
        nios_system_clock_5_out_read_last_time <= nios_system_clock_5_out_read;
    end


  //nios_system_clock_5_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_5_out_read != nios_system_clock_5_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_5_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_5_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_5_out_write_last_time <= 0;
      else 
        nios_system_clock_5_out_write_last_time <= nios_system_clock_5_out_write;
    end


  //nios_system_clock_5_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_5_out_write != nios_system_clock_5_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_5_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_5_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_5_out_writedata_last_time <= 0;
      else 
        nios_system_clock_5_out_writedata_last_time <= nios_system_clock_5_out_writedata;
    end


  //nios_system_clock_5_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_5_out_writedata != nios_system_clock_5_out_writedata_last_time) & nios_system_clock_5_out_write)
        begin
          $write("%0d ns: nios_system_clock_5_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_6_in_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_3_instruction_master_address_to_slave,
                                            cpu_3_instruction_master_dbs_address,
                                            cpu_3_instruction_master_latency_counter,
                                            cpu_3_instruction_master_read,
                                            cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                            nios_system_clock_6_in_endofpacket,
                                            nios_system_clock_6_in_readdata,
                                            nios_system_clock_6_in_waitrequest,
                                            reset_n,

                                           // outputs:
                                            cpu_3_instruction_master_granted_nios_system_clock_6_in,
                                            cpu_3_instruction_master_qualified_request_nios_system_clock_6_in,
                                            cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in,
                                            cpu_3_instruction_master_requests_nios_system_clock_6_in,
                                            d1_nios_system_clock_6_in_end_xfer,
                                            nios_system_clock_6_in_address,
                                            nios_system_clock_6_in_byteenable,
                                            nios_system_clock_6_in_endofpacket_from_sa,
                                            nios_system_clock_6_in_nativeaddress,
                                            nios_system_clock_6_in_read,
                                            nios_system_clock_6_in_readdata_from_sa,
                                            nios_system_clock_6_in_reset_n,
                                            nios_system_clock_6_in_waitrequest_from_sa,
                                            nios_system_clock_6_in_write
                                         )
;

  output           cpu_3_instruction_master_granted_nios_system_clock_6_in;
  output           cpu_3_instruction_master_qualified_request_nios_system_clock_6_in;
  output           cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in;
  output           cpu_3_instruction_master_requests_nios_system_clock_6_in;
  output           d1_nios_system_clock_6_in_end_xfer;
  output  [ 22: 0] nios_system_clock_6_in_address;
  output  [  1: 0] nios_system_clock_6_in_byteenable;
  output           nios_system_clock_6_in_endofpacket_from_sa;
  output  [ 21: 0] nios_system_clock_6_in_nativeaddress;
  output           nios_system_clock_6_in_read;
  output  [ 15: 0] nios_system_clock_6_in_readdata_from_sa;
  output           nios_system_clock_6_in_reset_n;
  output           nios_system_clock_6_in_waitrequest_from_sa;
  output           nios_system_clock_6_in_write;
  input            clk;
  input   [ 24: 0] cpu_3_instruction_master_address_to_slave;
  input   [  1: 0] cpu_3_instruction_master_dbs_address;
  input            cpu_3_instruction_master_latency_counter;
  input            cpu_3_instruction_master_read;
  input            cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            nios_system_clock_6_in_endofpacket;
  input   [ 15: 0] nios_system_clock_6_in_readdata;
  input            nios_system_clock_6_in_waitrequest;
  input            reset_n;

  wire             cpu_3_instruction_master_arbiterlock;
  wire             cpu_3_instruction_master_arbiterlock2;
  wire             cpu_3_instruction_master_continuerequest;
  wire             cpu_3_instruction_master_granted_nios_system_clock_6_in;
  wire             cpu_3_instruction_master_qualified_request_nios_system_clock_6_in;
  wire             cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in;
  wire             cpu_3_instruction_master_requests_nios_system_clock_6_in;
  wire             cpu_3_instruction_master_saved_grant_nios_system_clock_6_in;
  reg              d1_nios_system_clock_6_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_6_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 22: 0] nios_system_clock_6_in_address;
  wire             nios_system_clock_6_in_allgrants;
  wire             nios_system_clock_6_in_allow_new_arb_cycle;
  wire             nios_system_clock_6_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_6_in_any_continuerequest;
  wire             nios_system_clock_6_in_arb_counter_enable;
  reg     [  1: 0] nios_system_clock_6_in_arb_share_counter;
  wire    [  1: 0] nios_system_clock_6_in_arb_share_counter_next_value;
  wire    [  1: 0] nios_system_clock_6_in_arb_share_set_values;
  wire             nios_system_clock_6_in_beginbursttransfer_internal;
  wire             nios_system_clock_6_in_begins_xfer;
  wire    [  1: 0] nios_system_clock_6_in_byteenable;
  wire             nios_system_clock_6_in_end_xfer;
  wire             nios_system_clock_6_in_endofpacket_from_sa;
  wire             nios_system_clock_6_in_firsttransfer;
  wire             nios_system_clock_6_in_grant_vector;
  wire             nios_system_clock_6_in_in_a_read_cycle;
  wire             nios_system_clock_6_in_in_a_write_cycle;
  wire             nios_system_clock_6_in_master_qreq_vector;
  wire    [ 21: 0] nios_system_clock_6_in_nativeaddress;
  wire             nios_system_clock_6_in_non_bursting_master_requests;
  wire             nios_system_clock_6_in_read;
  wire    [ 15: 0] nios_system_clock_6_in_readdata_from_sa;
  reg              nios_system_clock_6_in_reg_firsttransfer;
  wire             nios_system_clock_6_in_reset_n;
  reg              nios_system_clock_6_in_slavearbiterlockenable;
  wire             nios_system_clock_6_in_slavearbiterlockenable2;
  wire             nios_system_clock_6_in_unreg_firsttransfer;
  wire             nios_system_clock_6_in_waitrequest_from_sa;
  wire             nios_system_clock_6_in_waits_for_read;
  wire             nios_system_clock_6_in_waits_for_write;
  wire             nios_system_clock_6_in_write;
  wire             wait_for_nios_system_clock_6_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_6_in_end_xfer;
    end


  assign nios_system_clock_6_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_3_instruction_master_qualified_request_nios_system_clock_6_in));
  //assign nios_system_clock_6_in_readdata_from_sa = nios_system_clock_6_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_6_in_readdata_from_sa = nios_system_clock_6_in_readdata;

  assign cpu_3_instruction_master_requests_nios_system_clock_6_in = (({cpu_3_instruction_master_address_to_slave[24 : 23] , 23'b0} == 25'h800000) & (cpu_3_instruction_master_read)) & cpu_3_instruction_master_read;
  //assign nios_system_clock_6_in_waitrequest_from_sa = nios_system_clock_6_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_6_in_waitrequest_from_sa = nios_system_clock_6_in_waitrequest;

  //nios_system_clock_6_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_6_in_arb_share_set_values = (cpu_3_instruction_master_granted_nios_system_clock_6_in)? 2 :
    1;

  //nios_system_clock_6_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_6_in_non_bursting_master_requests = cpu_3_instruction_master_requests_nios_system_clock_6_in;

  //nios_system_clock_6_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_6_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_6_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_6_in_arb_share_counter_next_value = nios_system_clock_6_in_firsttransfer ? (nios_system_clock_6_in_arb_share_set_values - 1) : |nios_system_clock_6_in_arb_share_counter ? (nios_system_clock_6_in_arb_share_counter - 1) : 0;

  //nios_system_clock_6_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_6_in_allgrants = |nios_system_clock_6_in_grant_vector;

  //nios_system_clock_6_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_6_in_end_xfer = ~(nios_system_clock_6_in_waits_for_read | nios_system_clock_6_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_6_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_6_in = nios_system_clock_6_in_end_xfer & (~nios_system_clock_6_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_6_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_6_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_6_in & nios_system_clock_6_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_6_in & ~nios_system_clock_6_in_non_bursting_master_requests);

  //nios_system_clock_6_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_6_in_arb_share_counter <= 0;
      else if (nios_system_clock_6_in_arb_counter_enable)
          nios_system_clock_6_in_arb_share_counter <= nios_system_clock_6_in_arb_share_counter_next_value;
    end


  //nios_system_clock_6_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_6_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_6_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_6_in) | (end_xfer_arb_share_counter_term_nios_system_clock_6_in & ~nios_system_clock_6_in_non_bursting_master_requests))
          nios_system_clock_6_in_slavearbiterlockenable <= |nios_system_clock_6_in_arb_share_counter_next_value;
    end


  //cpu_3/instruction_master nios_system_clock_6/in arbiterlock, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock = nios_system_clock_6_in_slavearbiterlockenable & cpu_3_instruction_master_continuerequest;

  //nios_system_clock_6_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_6_in_slavearbiterlockenable2 = |nios_system_clock_6_in_arb_share_counter_next_value;

  //cpu_3/instruction_master nios_system_clock_6/in arbiterlock2, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock2 = nios_system_clock_6_in_slavearbiterlockenable2 & cpu_3_instruction_master_continuerequest;

  //nios_system_clock_6_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_6_in_any_continuerequest = 1;

  //cpu_3_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_3_instruction_master_continuerequest = 1;

  assign cpu_3_instruction_master_qualified_request_nios_system_clock_6_in = cpu_3_instruction_master_requests_nios_system_clock_6_in & ~((cpu_3_instruction_master_read & ((cpu_3_instruction_master_latency_counter != 0) | (|cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))));
  //local readdatavalid cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in, which is an e_mux
  assign cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in = cpu_3_instruction_master_granted_nios_system_clock_6_in & cpu_3_instruction_master_read & ~nios_system_clock_6_in_waits_for_read;

  //assign nios_system_clock_6_in_endofpacket_from_sa = nios_system_clock_6_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_6_in_endofpacket_from_sa = nios_system_clock_6_in_endofpacket;

  //master is always granted when requested
  assign cpu_3_instruction_master_granted_nios_system_clock_6_in = cpu_3_instruction_master_qualified_request_nios_system_clock_6_in;

  //cpu_3/instruction_master saved-grant nios_system_clock_6/in, which is an e_assign
  assign cpu_3_instruction_master_saved_grant_nios_system_clock_6_in = cpu_3_instruction_master_requests_nios_system_clock_6_in;

  //allow new arb cycle for nios_system_clock_6/in, which is an e_assign
  assign nios_system_clock_6_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_6_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_6_in_master_qreq_vector = 1;

  //nios_system_clock_6_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_6_in_reset_n = reset_n;

  //nios_system_clock_6_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_6_in_firsttransfer = nios_system_clock_6_in_begins_xfer ? nios_system_clock_6_in_unreg_firsttransfer : nios_system_clock_6_in_reg_firsttransfer;

  //nios_system_clock_6_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_6_in_unreg_firsttransfer = ~(nios_system_clock_6_in_slavearbiterlockenable & nios_system_clock_6_in_any_continuerequest);

  //nios_system_clock_6_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_6_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_6_in_begins_xfer)
          nios_system_clock_6_in_reg_firsttransfer <= nios_system_clock_6_in_unreg_firsttransfer;
    end


  //nios_system_clock_6_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_6_in_beginbursttransfer_internal = nios_system_clock_6_in_begins_xfer;

  //nios_system_clock_6_in_read assignment, which is an e_mux
  assign nios_system_clock_6_in_read = cpu_3_instruction_master_granted_nios_system_clock_6_in & cpu_3_instruction_master_read;

  //nios_system_clock_6_in_write assignment, which is an e_mux
  assign nios_system_clock_6_in_write = 0;

  //nios_system_clock_6_in_address mux, which is an e_mux
  assign nios_system_clock_6_in_address = {cpu_3_instruction_master_address_to_slave >> 2,
    cpu_3_instruction_master_dbs_address[1],
    {1 {1'b0}}};

  //slaveid nios_system_clock_6_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_6_in_nativeaddress = cpu_3_instruction_master_address_to_slave >> 2;

  //d1_nios_system_clock_6_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_6_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_6_in_end_xfer <= nios_system_clock_6_in_end_xfer;
    end


  //nios_system_clock_6_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_6_in_waits_for_read = nios_system_clock_6_in_in_a_read_cycle & nios_system_clock_6_in_waitrequest_from_sa;

  //nios_system_clock_6_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_6_in_in_a_read_cycle = cpu_3_instruction_master_granted_nios_system_clock_6_in & cpu_3_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_6_in_in_a_read_cycle;

  //nios_system_clock_6_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_6_in_waits_for_write = nios_system_clock_6_in_in_a_write_cycle & nios_system_clock_6_in_waitrequest_from_sa;

  //nios_system_clock_6_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_6_in_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_6_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_6_in_counter = 0;
  //nios_system_clock_6_in_byteenable byte enable port mux, which is an e_mux
  assign nios_system_clock_6_in_byteenable = -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_6/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_6_out_arbitrator (
                                            // inputs:
                                             clk,
                                             d1_sdram_0_s1_end_xfer,
                                             nios_system_clock_6_out_address,
                                             nios_system_clock_6_out_byteenable,
                                             nios_system_clock_6_out_granted_sdram_0_s1,
                                             nios_system_clock_6_out_qualified_request_sdram_0_s1,
                                             nios_system_clock_6_out_read,
                                             nios_system_clock_6_out_read_data_valid_sdram_0_s1,
                                             nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register,
                                             nios_system_clock_6_out_requests_sdram_0_s1,
                                             nios_system_clock_6_out_write,
                                             nios_system_clock_6_out_writedata,
                                             reset_n,
                                             sdram_0_s1_readdata_from_sa,
                                             sdram_0_s1_waitrequest_from_sa,

                                            // outputs:
                                             nios_system_clock_6_out_address_to_slave,
                                             nios_system_clock_6_out_readdata,
                                             nios_system_clock_6_out_reset_n,
                                             nios_system_clock_6_out_waitrequest
                                          )
;

  output  [ 22: 0] nios_system_clock_6_out_address_to_slave;
  output  [ 15: 0] nios_system_clock_6_out_readdata;
  output           nios_system_clock_6_out_reset_n;
  output           nios_system_clock_6_out_waitrequest;
  input            clk;
  input            d1_sdram_0_s1_end_xfer;
  input   [ 22: 0] nios_system_clock_6_out_address;
  input   [  1: 0] nios_system_clock_6_out_byteenable;
  input            nios_system_clock_6_out_granted_sdram_0_s1;
  input            nios_system_clock_6_out_qualified_request_sdram_0_s1;
  input            nios_system_clock_6_out_read;
  input            nios_system_clock_6_out_read_data_valid_sdram_0_s1;
  input            nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register;
  input            nios_system_clock_6_out_requests_sdram_0_s1;
  input            nios_system_clock_6_out_write;
  input   [ 15: 0] nios_system_clock_6_out_writedata;
  input            reset_n;
  input   [ 15: 0] sdram_0_s1_readdata_from_sa;
  input            sdram_0_s1_waitrequest_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 22: 0] nios_system_clock_6_out_address_last_time;
  wire    [ 22: 0] nios_system_clock_6_out_address_to_slave;
  reg     [  1: 0] nios_system_clock_6_out_byteenable_last_time;
  reg              nios_system_clock_6_out_read_last_time;
  wire    [ 15: 0] nios_system_clock_6_out_readdata;
  wire             nios_system_clock_6_out_reset_n;
  wire             nios_system_clock_6_out_run;
  wire             nios_system_clock_6_out_waitrequest;
  reg              nios_system_clock_6_out_write_last_time;
  reg     [ 15: 0] nios_system_clock_6_out_writedata_last_time;
  wire             r_3;
  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (nios_system_clock_6_out_qualified_request_sdram_0_s1 | nios_system_clock_6_out_read_data_valid_sdram_0_s1 | ~nios_system_clock_6_out_requests_sdram_0_s1) & (nios_system_clock_6_out_granted_sdram_0_s1 | ~nios_system_clock_6_out_qualified_request_sdram_0_s1) & ((~nios_system_clock_6_out_qualified_request_sdram_0_s1 | ~nios_system_clock_6_out_read | (nios_system_clock_6_out_read_data_valid_sdram_0_s1 & nios_system_clock_6_out_read))) & ((~nios_system_clock_6_out_qualified_request_sdram_0_s1 | ~(nios_system_clock_6_out_read | nios_system_clock_6_out_write) | (1 & ~sdram_0_s1_waitrequest_from_sa & (nios_system_clock_6_out_read | nios_system_clock_6_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_6_out_run = r_3;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_6_out_address_to_slave = nios_system_clock_6_out_address;

  //nios_system_clock_6/out readdata mux, which is an e_mux
  assign nios_system_clock_6_out_readdata = sdram_0_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_6_out_waitrequest = ~nios_system_clock_6_out_run;

  //nios_system_clock_6_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_6_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_6_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_6_out_address_last_time <= 0;
      else 
        nios_system_clock_6_out_address_last_time <= nios_system_clock_6_out_address;
    end


  //nios_system_clock_6/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_6_out_waitrequest & (nios_system_clock_6_out_read | nios_system_clock_6_out_write);
    end


  //nios_system_clock_6_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_6_out_address != nios_system_clock_6_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_6_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_6_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_6_out_byteenable_last_time <= 0;
      else 
        nios_system_clock_6_out_byteenable_last_time <= nios_system_clock_6_out_byteenable;
    end


  //nios_system_clock_6_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_6_out_byteenable != nios_system_clock_6_out_byteenable_last_time))
        begin
          $write("%0d ns: nios_system_clock_6_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_6_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_6_out_read_last_time <= 0;
      else 
        nios_system_clock_6_out_read_last_time <= nios_system_clock_6_out_read;
    end


  //nios_system_clock_6_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_6_out_read != nios_system_clock_6_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_6_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_6_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_6_out_write_last_time <= 0;
      else 
        nios_system_clock_6_out_write_last_time <= nios_system_clock_6_out_write;
    end


  //nios_system_clock_6_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_6_out_write != nios_system_clock_6_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_6_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_6_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_6_out_writedata_last_time <= 0;
      else 
        nios_system_clock_6_out_writedata_last_time <= nios_system_clock_6_out_writedata;
    end


  //nios_system_clock_6_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_6_out_writedata != nios_system_clock_6_out_writedata_last_time) & nios_system_clock_6_out_write)
        begin
          $write("%0d ns: nios_system_clock_6_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_7_in_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_3_data_master_address_to_slave,
                                            cpu_3_data_master_byteenable,
                                            cpu_3_data_master_dbs_address,
                                            cpu_3_data_master_dbs_write_16,
                                            cpu_3_data_master_latency_counter,
                                            cpu_3_data_master_read,
                                            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                            cpu_3_data_master_write,
                                            nios_system_clock_7_in_endofpacket,
                                            nios_system_clock_7_in_readdata,
                                            nios_system_clock_7_in_waitrequest,
                                            reset_n,

                                           // outputs:
                                            cpu_3_data_master_byteenable_nios_system_clock_7_in,
                                            cpu_3_data_master_granted_nios_system_clock_7_in,
                                            cpu_3_data_master_qualified_request_nios_system_clock_7_in,
                                            cpu_3_data_master_read_data_valid_nios_system_clock_7_in,
                                            cpu_3_data_master_requests_nios_system_clock_7_in,
                                            d1_nios_system_clock_7_in_end_xfer,
                                            nios_system_clock_7_in_address,
                                            nios_system_clock_7_in_byteenable,
                                            nios_system_clock_7_in_endofpacket_from_sa,
                                            nios_system_clock_7_in_nativeaddress,
                                            nios_system_clock_7_in_read,
                                            nios_system_clock_7_in_readdata_from_sa,
                                            nios_system_clock_7_in_reset_n,
                                            nios_system_clock_7_in_waitrequest_from_sa,
                                            nios_system_clock_7_in_write,
                                            nios_system_clock_7_in_writedata
                                         )
;

  output  [  1: 0] cpu_3_data_master_byteenable_nios_system_clock_7_in;
  output           cpu_3_data_master_granted_nios_system_clock_7_in;
  output           cpu_3_data_master_qualified_request_nios_system_clock_7_in;
  output           cpu_3_data_master_read_data_valid_nios_system_clock_7_in;
  output           cpu_3_data_master_requests_nios_system_clock_7_in;
  output           d1_nios_system_clock_7_in_end_xfer;
  output  [ 22: 0] nios_system_clock_7_in_address;
  output  [  1: 0] nios_system_clock_7_in_byteenable;
  output           nios_system_clock_7_in_endofpacket_from_sa;
  output  [ 21: 0] nios_system_clock_7_in_nativeaddress;
  output           nios_system_clock_7_in_read;
  output  [ 15: 0] nios_system_clock_7_in_readdata_from_sa;
  output           nios_system_clock_7_in_reset_n;
  output           nios_system_clock_7_in_waitrequest_from_sa;
  output           nios_system_clock_7_in_write;
  output  [ 15: 0] nios_system_clock_7_in_writedata;
  input            clk;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input   [  3: 0] cpu_3_data_master_byteenable;
  input   [  1: 0] cpu_3_data_master_dbs_address;
  input   [ 15: 0] cpu_3_data_master_dbs_write_16;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input            nios_system_clock_7_in_endofpacket;
  input   [ 15: 0] nios_system_clock_7_in_readdata;
  input            nios_system_clock_7_in_waitrequest;
  input            reset_n;

  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire    [  1: 0] cpu_3_data_master_byteenable_nios_system_clock_7_in;
  wire    [  1: 0] cpu_3_data_master_byteenable_nios_system_clock_7_in_segment_0;
  wire    [  1: 0] cpu_3_data_master_byteenable_nios_system_clock_7_in_segment_1;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_nios_system_clock_7_in;
  wire             cpu_3_data_master_qualified_request_nios_system_clock_7_in;
  wire             cpu_3_data_master_read_data_valid_nios_system_clock_7_in;
  wire             cpu_3_data_master_requests_nios_system_clock_7_in;
  wire             cpu_3_data_master_saved_grant_nios_system_clock_7_in;
  reg              d1_nios_system_clock_7_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_7_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 22: 0] nios_system_clock_7_in_address;
  wire             nios_system_clock_7_in_allgrants;
  wire             nios_system_clock_7_in_allow_new_arb_cycle;
  wire             nios_system_clock_7_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_7_in_any_continuerequest;
  wire             nios_system_clock_7_in_arb_counter_enable;
  reg     [  2: 0] nios_system_clock_7_in_arb_share_counter;
  wire    [  2: 0] nios_system_clock_7_in_arb_share_counter_next_value;
  wire    [  2: 0] nios_system_clock_7_in_arb_share_set_values;
  wire             nios_system_clock_7_in_beginbursttransfer_internal;
  wire             nios_system_clock_7_in_begins_xfer;
  wire    [  1: 0] nios_system_clock_7_in_byteenable;
  wire             nios_system_clock_7_in_end_xfer;
  wire             nios_system_clock_7_in_endofpacket_from_sa;
  wire             nios_system_clock_7_in_firsttransfer;
  wire             nios_system_clock_7_in_grant_vector;
  wire             nios_system_clock_7_in_in_a_read_cycle;
  wire             nios_system_clock_7_in_in_a_write_cycle;
  wire             nios_system_clock_7_in_master_qreq_vector;
  wire    [ 21: 0] nios_system_clock_7_in_nativeaddress;
  wire             nios_system_clock_7_in_non_bursting_master_requests;
  wire             nios_system_clock_7_in_read;
  wire    [ 15: 0] nios_system_clock_7_in_readdata_from_sa;
  reg              nios_system_clock_7_in_reg_firsttransfer;
  wire             nios_system_clock_7_in_reset_n;
  reg              nios_system_clock_7_in_slavearbiterlockenable;
  wire             nios_system_clock_7_in_slavearbiterlockenable2;
  wire             nios_system_clock_7_in_unreg_firsttransfer;
  wire             nios_system_clock_7_in_waitrequest_from_sa;
  wire             nios_system_clock_7_in_waits_for_read;
  wire             nios_system_clock_7_in_waits_for_write;
  wire             nios_system_clock_7_in_write;
  wire    [ 15: 0] nios_system_clock_7_in_writedata;
  wire             wait_for_nios_system_clock_7_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_7_in_end_xfer;
    end


  assign nios_system_clock_7_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_3_data_master_qualified_request_nios_system_clock_7_in));
  //assign nios_system_clock_7_in_readdata_from_sa = nios_system_clock_7_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_7_in_readdata_from_sa = nios_system_clock_7_in_readdata;

  assign cpu_3_data_master_requests_nios_system_clock_7_in = ({cpu_3_data_master_address_to_slave[24 : 23] , 23'b0} == 25'h800000) & (cpu_3_data_master_read | cpu_3_data_master_write);
  //assign nios_system_clock_7_in_waitrequest_from_sa = nios_system_clock_7_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_7_in_waitrequest_from_sa = nios_system_clock_7_in_waitrequest;

  //nios_system_clock_7_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_7_in_arb_share_set_values = (cpu_3_data_master_granted_nios_system_clock_7_in)? 2 :
    1;

  //nios_system_clock_7_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_7_in_non_bursting_master_requests = cpu_3_data_master_requests_nios_system_clock_7_in;

  //nios_system_clock_7_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_7_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_7_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_7_in_arb_share_counter_next_value = nios_system_clock_7_in_firsttransfer ? (nios_system_clock_7_in_arb_share_set_values - 1) : |nios_system_clock_7_in_arb_share_counter ? (nios_system_clock_7_in_arb_share_counter - 1) : 0;

  //nios_system_clock_7_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_7_in_allgrants = |nios_system_clock_7_in_grant_vector;

  //nios_system_clock_7_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_7_in_end_xfer = ~(nios_system_clock_7_in_waits_for_read | nios_system_clock_7_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_7_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_7_in = nios_system_clock_7_in_end_xfer & (~nios_system_clock_7_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_7_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_7_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_7_in & nios_system_clock_7_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_7_in & ~nios_system_clock_7_in_non_bursting_master_requests);

  //nios_system_clock_7_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_7_in_arb_share_counter <= 0;
      else if (nios_system_clock_7_in_arb_counter_enable)
          nios_system_clock_7_in_arb_share_counter <= nios_system_clock_7_in_arb_share_counter_next_value;
    end


  //nios_system_clock_7_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_7_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_7_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_7_in) | (end_xfer_arb_share_counter_term_nios_system_clock_7_in & ~nios_system_clock_7_in_non_bursting_master_requests))
          nios_system_clock_7_in_slavearbiterlockenable <= |nios_system_clock_7_in_arb_share_counter_next_value;
    end


  //cpu_3/data_master nios_system_clock_7/in arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = nios_system_clock_7_in_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //nios_system_clock_7_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_7_in_slavearbiterlockenable2 = |nios_system_clock_7_in_arb_share_counter_next_value;

  //cpu_3/data_master nios_system_clock_7/in arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = nios_system_clock_7_in_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //nios_system_clock_7_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_7_in_any_continuerequest = 1;

  //cpu_3_data_master_continuerequest continued request, which is an e_assign
  assign cpu_3_data_master_continuerequest = 1;

  assign cpu_3_data_master_qualified_request_nios_system_clock_7_in = cpu_3_data_master_requests_nios_system_clock_7_in & ~((cpu_3_data_master_read & ((cpu_3_data_master_latency_counter != 0) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | ((!cpu_3_data_master_byteenable_nios_system_clock_7_in) & cpu_3_data_master_write));
  //local readdatavalid cpu_3_data_master_read_data_valid_nios_system_clock_7_in, which is an e_mux
  assign cpu_3_data_master_read_data_valid_nios_system_clock_7_in = cpu_3_data_master_granted_nios_system_clock_7_in & cpu_3_data_master_read & ~nios_system_clock_7_in_waits_for_read;

  //nios_system_clock_7_in_writedata mux, which is an e_mux
  assign nios_system_clock_7_in_writedata = cpu_3_data_master_dbs_write_16;

  //assign nios_system_clock_7_in_endofpacket_from_sa = nios_system_clock_7_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_7_in_endofpacket_from_sa = nios_system_clock_7_in_endofpacket;

  //master is always granted when requested
  assign cpu_3_data_master_granted_nios_system_clock_7_in = cpu_3_data_master_qualified_request_nios_system_clock_7_in;

  //cpu_3/data_master saved-grant nios_system_clock_7/in, which is an e_assign
  assign cpu_3_data_master_saved_grant_nios_system_clock_7_in = cpu_3_data_master_requests_nios_system_clock_7_in;

  //allow new arb cycle for nios_system_clock_7/in, which is an e_assign
  assign nios_system_clock_7_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_7_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_7_in_master_qreq_vector = 1;

  //nios_system_clock_7_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_7_in_reset_n = reset_n;

  //nios_system_clock_7_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_7_in_firsttransfer = nios_system_clock_7_in_begins_xfer ? nios_system_clock_7_in_unreg_firsttransfer : nios_system_clock_7_in_reg_firsttransfer;

  //nios_system_clock_7_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_7_in_unreg_firsttransfer = ~(nios_system_clock_7_in_slavearbiterlockenable & nios_system_clock_7_in_any_continuerequest);

  //nios_system_clock_7_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_7_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_7_in_begins_xfer)
          nios_system_clock_7_in_reg_firsttransfer <= nios_system_clock_7_in_unreg_firsttransfer;
    end


  //nios_system_clock_7_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_7_in_beginbursttransfer_internal = nios_system_clock_7_in_begins_xfer;

  //nios_system_clock_7_in_read assignment, which is an e_mux
  assign nios_system_clock_7_in_read = cpu_3_data_master_granted_nios_system_clock_7_in & cpu_3_data_master_read;

  //nios_system_clock_7_in_write assignment, which is an e_mux
  assign nios_system_clock_7_in_write = cpu_3_data_master_granted_nios_system_clock_7_in & cpu_3_data_master_write;

  //nios_system_clock_7_in_address mux, which is an e_mux
  assign nios_system_clock_7_in_address = {cpu_3_data_master_address_to_slave >> 2,
    cpu_3_data_master_dbs_address[1],
    {1 {1'b0}}};

  //slaveid nios_system_clock_7_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_7_in_nativeaddress = cpu_3_data_master_address_to_slave >> 2;

  //d1_nios_system_clock_7_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_7_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_7_in_end_xfer <= nios_system_clock_7_in_end_xfer;
    end


  //nios_system_clock_7_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_7_in_waits_for_read = nios_system_clock_7_in_in_a_read_cycle & nios_system_clock_7_in_waitrequest_from_sa;

  //nios_system_clock_7_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_7_in_in_a_read_cycle = cpu_3_data_master_granted_nios_system_clock_7_in & cpu_3_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_7_in_in_a_read_cycle;

  //nios_system_clock_7_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_7_in_waits_for_write = nios_system_clock_7_in_in_a_write_cycle & nios_system_clock_7_in_waitrequest_from_sa;

  //nios_system_clock_7_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_7_in_in_a_write_cycle = cpu_3_data_master_granted_nios_system_clock_7_in & cpu_3_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_7_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_7_in_counter = 0;
  //nios_system_clock_7_in_byteenable byte enable port mux, which is an e_mux
  assign nios_system_clock_7_in_byteenable = (cpu_3_data_master_granted_nios_system_clock_7_in)? cpu_3_data_master_byteenable_nios_system_clock_7_in :
    -1;

  assign {cpu_3_data_master_byteenable_nios_system_clock_7_in_segment_1,
cpu_3_data_master_byteenable_nios_system_clock_7_in_segment_0} = cpu_3_data_master_byteenable;
  assign cpu_3_data_master_byteenable_nios_system_clock_7_in = ((cpu_3_data_master_dbs_address[1] == 0))? cpu_3_data_master_byteenable_nios_system_clock_7_in_segment_0 :
    cpu_3_data_master_byteenable_nios_system_clock_7_in_segment_1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_7/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_7_out_arbitrator (
                                            // inputs:
                                             clk,
                                             d1_sdram_0_s1_end_xfer,
                                             nios_system_clock_7_out_address,
                                             nios_system_clock_7_out_byteenable,
                                             nios_system_clock_7_out_granted_sdram_0_s1,
                                             nios_system_clock_7_out_qualified_request_sdram_0_s1,
                                             nios_system_clock_7_out_read,
                                             nios_system_clock_7_out_read_data_valid_sdram_0_s1,
                                             nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register,
                                             nios_system_clock_7_out_requests_sdram_0_s1,
                                             nios_system_clock_7_out_write,
                                             nios_system_clock_7_out_writedata,
                                             reset_n,
                                             sdram_0_s1_readdata_from_sa,
                                             sdram_0_s1_waitrequest_from_sa,

                                            // outputs:
                                             nios_system_clock_7_out_address_to_slave,
                                             nios_system_clock_7_out_readdata,
                                             nios_system_clock_7_out_reset_n,
                                             nios_system_clock_7_out_waitrequest
                                          )
;

  output  [ 22: 0] nios_system_clock_7_out_address_to_slave;
  output  [ 15: 0] nios_system_clock_7_out_readdata;
  output           nios_system_clock_7_out_reset_n;
  output           nios_system_clock_7_out_waitrequest;
  input            clk;
  input            d1_sdram_0_s1_end_xfer;
  input   [ 22: 0] nios_system_clock_7_out_address;
  input   [  1: 0] nios_system_clock_7_out_byteenable;
  input            nios_system_clock_7_out_granted_sdram_0_s1;
  input            nios_system_clock_7_out_qualified_request_sdram_0_s1;
  input            nios_system_clock_7_out_read;
  input            nios_system_clock_7_out_read_data_valid_sdram_0_s1;
  input            nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register;
  input            nios_system_clock_7_out_requests_sdram_0_s1;
  input            nios_system_clock_7_out_write;
  input   [ 15: 0] nios_system_clock_7_out_writedata;
  input            reset_n;
  input   [ 15: 0] sdram_0_s1_readdata_from_sa;
  input            sdram_0_s1_waitrequest_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 22: 0] nios_system_clock_7_out_address_last_time;
  wire    [ 22: 0] nios_system_clock_7_out_address_to_slave;
  reg     [  1: 0] nios_system_clock_7_out_byteenable_last_time;
  reg              nios_system_clock_7_out_read_last_time;
  wire    [ 15: 0] nios_system_clock_7_out_readdata;
  wire             nios_system_clock_7_out_reset_n;
  wire             nios_system_clock_7_out_run;
  wire             nios_system_clock_7_out_waitrequest;
  reg              nios_system_clock_7_out_write_last_time;
  reg     [ 15: 0] nios_system_clock_7_out_writedata_last_time;
  wire             r_3;
  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (nios_system_clock_7_out_qualified_request_sdram_0_s1 | nios_system_clock_7_out_read_data_valid_sdram_0_s1 | ~nios_system_clock_7_out_requests_sdram_0_s1) & (nios_system_clock_7_out_granted_sdram_0_s1 | ~nios_system_clock_7_out_qualified_request_sdram_0_s1) & ((~nios_system_clock_7_out_qualified_request_sdram_0_s1 | ~nios_system_clock_7_out_read | (nios_system_clock_7_out_read_data_valid_sdram_0_s1 & nios_system_clock_7_out_read))) & ((~nios_system_clock_7_out_qualified_request_sdram_0_s1 | ~(nios_system_clock_7_out_read | nios_system_clock_7_out_write) | (1 & ~sdram_0_s1_waitrequest_from_sa & (nios_system_clock_7_out_read | nios_system_clock_7_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_7_out_run = r_3;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_7_out_address_to_slave = nios_system_clock_7_out_address;

  //nios_system_clock_7/out readdata mux, which is an e_mux
  assign nios_system_clock_7_out_readdata = sdram_0_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_7_out_waitrequest = ~nios_system_clock_7_out_run;

  //nios_system_clock_7_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_7_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_7_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_7_out_address_last_time <= 0;
      else 
        nios_system_clock_7_out_address_last_time <= nios_system_clock_7_out_address;
    end


  //nios_system_clock_7/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_7_out_waitrequest & (nios_system_clock_7_out_read | nios_system_clock_7_out_write);
    end


  //nios_system_clock_7_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_7_out_address != nios_system_clock_7_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_7_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_7_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_7_out_byteenable_last_time <= 0;
      else 
        nios_system_clock_7_out_byteenable_last_time <= nios_system_clock_7_out_byteenable;
    end


  //nios_system_clock_7_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_7_out_byteenable != nios_system_clock_7_out_byteenable_last_time))
        begin
          $write("%0d ns: nios_system_clock_7_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_7_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_7_out_read_last_time <= 0;
      else 
        nios_system_clock_7_out_read_last_time <= nios_system_clock_7_out_read;
    end


  //nios_system_clock_7_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_7_out_read != nios_system_clock_7_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_7_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_7_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_7_out_write_last_time <= 0;
      else 
        nios_system_clock_7_out_write_last_time <= nios_system_clock_7_out_write;
    end


  //nios_system_clock_7_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_7_out_write != nios_system_clock_7_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_7_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_7_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_7_out_writedata_last_time <= 0;
      else 
        nios_system_clock_7_out_writedata_last_time <= nios_system_clock_7_out_writedata;
    end


  //nios_system_clock_7_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_7_out_writedata != nios_system_clock_7_out_writedata_last_time) & nios_system_clock_7_out_write)
        begin
          $write("%0d ns: nios_system_clock_7_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_8_in_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_1_data_master_address_to_slave,
                                            cpu_1_data_master_byteenable,
                                            cpu_1_data_master_dbs_address,
                                            cpu_1_data_master_dbs_write_8,
                                            cpu_1_data_master_latency_counter,
                                            cpu_1_data_master_read,
                                            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                            cpu_1_data_master_write,
                                            nios_system_clock_8_in_endofpacket,
                                            nios_system_clock_8_in_readdata,
                                            nios_system_clock_8_in_waitrequest,
                                            reset_n,

                                           // outputs:
                                            cpu_1_data_master_byteenable_nios_system_clock_8_in,
                                            cpu_1_data_master_granted_nios_system_clock_8_in,
                                            cpu_1_data_master_qualified_request_nios_system_clock_8_in,
                                            cpu_1_data_master_read_data_valid_nios_system_clock_8_in,
                                            cpu_1_data_master_requests_nios_system_clock_8_in,
                                            d1_nios_system_clock_8_in_end_xfer,
                                            nios_system_clock_8_in_address,
                                            nios_system_clock_8_in_endofpacket_from_sa,
                                            nios_system_clock_8_in_nativeaddress,
                                            nios_system_clock_8_in_read,
                                            nios_system_clock_8_in_readdata_from_sa,
                                            nios_system_clock_8_in_reset_n,
                                            nios_system_clock_8_in_waitrequest_from_sa,
                                            nios_system_clock_8_in_write,
                                            nios_system_clock_8_in_writedata
                                         )
;

  output           cpu_1_data_master_byteenable_nios_system_clock_8_in;
  output           cpu_1_data_master_granted_nios_system_clock_8_in;
  output           cpu_1_data_master_qualified_request_nios_system_clock_8_in;
  output           cpu_1_data_master_read_data_valid_nios_system_clock_8_in;
  output           cpu_1_data_master_requests_nios_system_clock_8_in;
  output           d1_nios_system_clock_8_in_end_xfer;
  output           nios_system_clock_8_in_address;
  output           nios_system_clock_8_in_endofpacket_from_sa;
  output           nios_system_clock_8_in_nativeaddress;
  output           nios_system_clock_8_in_read;
  output  [  7: 0] nios_system_clock_8_in_readdata_from_sa;
  output           nios_system_clock_8_in_reset_n;
  output           nios_system_clock_8_in_waitrequest_from_sa;
  output           nios_system_clock_8_in_write;
  output  [  7: 0] nios_system_clock_8_in_writedata;
  input            clk;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input   [  3: 0] cpu_1_data_master_byteenable;
  input   [  1: 0] cpu_1_data_master_dbs_address;
  input   [  7: 0] cpu_1_data_master_dbs_write_8;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input            nios_system_clock_8_in_endofpacket;
  input   [  7: 0] nios_system_clock_8_in_readdata;
  input            nios_system_clock_8_in_waitrequest;
  input            reset_n;

  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_byteenable_nios_system_clock_8_in;
  wire             cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_0;
  wire             cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_1;
  wire             cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_2;
  wire             cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_3;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_nios_system_clock_8_in;
  wire             cpu_1_data_master_qualified_request_nios_system_clock_8_in;
  wire             cpu_1_data_master_read_data_valid_nios_system_clock_8_in;
  wire             cpu_1_data_master_requests_nios_system_clock_8_in;
  wire             cpu_1_data_master_saved_grant_nios_system_clock_8_in;
  reg              d1_nios_system_clock_8_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_8_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             nios_system_clock_8_in_address;
  wire             nios_system_clock_8_in_allgrants;
  wire             nios_system_clock_8_in_allow_new_arb_cycle;
  wire             nios_system_clock_8_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_8_in_any_continuerequest;
  wire             nios_system_clock_8_in_arb_counter_enable;
  reg     [  2: 0] nios_system_clock_8_in_arb_share_counter;
  wire    [  2: 0] nios_system_clock_8_in_arb_share_counter_next_value;
  wire    [  2: 0] nios_system_clock_8_in_arb_share_set_values;
  wire             nios_system_clock_8_in_beginbursttransfer_internal;
  wire             nios_system_clock_8_in_begins_xfer;
  wire             nios_system_clock_8_in_end_xfer;
  wire             nios_system_clock_8_in_endofpacket_from_sa;
  wire             nios_system_clock_8_in_firsttransfer;
  wire             nios_system_clock_8_in_grant_vector;
  wire             nios_system_clock_8_in_in_a_read_cycle;
  wire             nios_system_clock_8_in_in_a_write_cycle;
  wire             nios_system_clock_8_in_master_qreq_vector;
  wire             nios_system_clock_8_in_nativeaddress;
  wire             nios_system_clock_8_in_non_bursting_master_requests;
  wire             nios_system_clock_8_in_pretend_byte_enable;
  wire             nios_system_clock_8_in_read;
  wire    [  7: 0] nios_system_clock_8_in_readdata_from_sa;
  reg              nios_system_clock_8_in_reg_firsttransfer;
  wire             nios_system_clock_8_in_reset_n;
  reg              nios_system_clock_8_in_slavearbiterlockenable;
  wire             nios_system_clock_8_in_slavearbiterlockenable2;
  wire             nios_system_clock_8_in_unreg_firsttransfer;
  wire             nios_system_clock_8_in_waitrequest_from_sa;
  wire             nios_system_clock_8_in_waits_for_read;
  wire             nios_system_clock_8_in_waits_for_write;
  wire             nios_system_clock_8_in_write;
  wire    [  7: 0] nios_system_clock_8_in_writedata;
  wire             wait_for_nios_system_clock_8_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_8_in_end_xfer;
    end


  assign nios_system_clock_8_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_1_data_master_qualified_request_nios_system_clock_8_in));
  //assign nios_system_clock_8_in_readdata_from_sa = nios_system_clock_8_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_8_in_readdata_from_sa = nios_system_clock_8_in_readdata;

  assign cpu_1_data_master_requests_nios_system_clock_8_in = ({cpu_1_data_master_address_to_slave[24 : 1] , 1'b0} == 25'h19030d8) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //assign nios_system_clock_8_in_waitrequest_from_sa = nios_system_clock_8_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_8_in_waitrequest_from_sa = nios_system_clock_8_in_waitrequest;

  //nios_system_clock_8_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_8_in_arb_share_set_values = (cpu_1_data_master_granted_nios_system_clock_8_in)? 4 :
    1;

  //nios_system_clock_8_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_8_in_non_bursting_master_requests = cpu_1_data_master_requests_nios_system_clock_8_in;

  //nios_system_clock_8_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_8_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_8_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_8_in_arb_share_counter_next_value = nios_system_clock_8_in_firsttransfer ? (nios_system_clock_8_in_arb_share_set_values - 1) : |nios_system_clock_8_in_arb_share_counter ? (nios_system_clock_8_in_arb_share_counter - 1) : 0;

  //nios_system_clock_8_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_8_in_allgrants = |nios_system_clock_8_in_grant_vector;

  //nios_system_clock_8_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_8_in_end_xfer = ~(nios_system_clock_8_in_waits_for_read | nios_system_clock_8_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_8_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_8_in = nios_system_clock_8_in_end_xfer & (~nios_system_clock_8_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_8_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_8_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_8_in & nios_system_clock_8_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_8_in & ~nios_system_clock_8_in_non_bursting_master_requests);

  //nios_system_clock_8_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_8_in_arb_share_counter <= 0;
      else if (nios_system_clock_8_in_arb_counter_enable)
          nios_system_clock_8_in_arb_share_counter <= nios_system_clock_8_in_arb_share_counter_next_value;
    end


  //nios_system_clock_8_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_8_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_8_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_8_in) | (end_xfer_arb_share_counter_term_nios_system_clock_8_in & ~nios_system_clock_8_in_non_bursting_master_requests))
          nios_system_clock_8_in_slavearbiterlockenable <= |nios_system_clock_8_in_arb_share_counter_next_value;
    end


  //cpu_1/data_master nios_system_clock_8/in arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = nios_system_clock_8_in_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //nios_system_clock_8_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_8_in_slavearbiterlockenable2 = |nios_system_clock_8_in_arb_share_counter_next_value;

  //cpu_1/data_master nios_system_clock_8/in arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = nios_system_clock_8_in_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //nios_system_clock_8_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_8_in_any_continuerequest = 1;

  //cpu_1_data_master_continuerequest continued request, which is an e_assign
  assign cpu_1_data_master_continuerequest = 1;

  assign cpu_1_data_master_qualified_request_nios_system_clock_8_in = cpu_1_data_master_requests_nios_system_clock_8_in & ~((cpu_1_data_master_read & ((cpu_1_data_master_latency_counter != 0) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | ((!cpu_1_data_master_byteenable_nios_system_clock_8_in) & cpu_1_data_master_write));
  //local readdatavalid cpu_1_data_master_read_data_valid_nios_system_clock_8_in, which is an e_mux
  assign cpu_1_data_master_read_data_valid_nios_system_clock_8_in = cpu_1_data_master_granted_nios_system_clock_8_in & cpu_1_data_master_read & ~nios_system_clock_8_in_waits_for_read;

  //nios_system_clock_8_in_writedata mux, which is an e_mux
  assign nios_system_clock_8_in_writedata = cpu_1_data_master_dbs_write_8;

  //assign nios_system_clock_8_in_endofpacket_from_sa = nios_system_clock_8_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_8_in_endofpacket_from_sa = nios_system_clock_8_in_endofpacket;

  //master is always granted when requested
  assign cpu_1_data_master_granted_nios_system_clock_8_in = cpu_1_data_master_qualified_request_nios_system_clock_8_in;

  //cpu_1/data_master saved-grant nios_system_clock_8/in, which is an e_assign
  assign cpu_1_data_master_saved_grant_nios_system_clock_8_in = cpu_1_data_master_requests_nios_system_clock_8_in;

  //allow new arb cycle for nios_system_clock_8/in, which is an e_assign
  assign nios_system_clock_8_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_8_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_8_in_master_qreq_vector = 1;

  //nios_system_clock_8_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_8_in_reset_n = reset_n;

  //nios_system_clock_8_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_8_in_firsttransfer = nios_system_clock_8_in_begins_xfer ? nios_system_clock_8_in_unreg_firsttransfer : nios_system_clock_8_in_reg_firsttransfer;

  //nios_system_clock_8_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_8_in_unreg_firsttransfer = ~(nios_system_clock_8_in_slavearbiterlockenable & nios_system_clock_8_in_any_continuerequest);

  //nios_system_clock_8_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_8_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_8_in_begins_xfer)
          nios_system_clock_8_in_reg_firsttransfer <= nios_system_clock_8_in_unreg_firsttransfer;
    end


  //nios_system_clock_8_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_8_in_beginbursttransfer_internal = nios_system_clock_8_in_begins_xfer;

  //nios_system_clock_8_in_read assignment, which is an e_mux
  assign nios_system_clock_8_in_read = cpu_1_data_master_granted_nios_system_clock_8_in & cpu_1_data_master_read;

  //nios_system_clock_8_in_write assignment, which is an e_mux
  assign nios_system_clock_8_in_write = ((cpu_1_data_master_granted_nios_system_clock_8_in & cpu_1_data_master_write)) & nios_system_clock_8_in_pretend_byte_enable;

  //nios_system_clock_8_in_address mux, which is an e_mux
  assign nios_system_clock_8_in_address = {cpu_1_data_master_address_to_slave >> 2,
    cpu_1_data_master_dbs_address[1 : 0]};

  //slaveid nios_system_clock_8_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_8_in_nativeaddress = cpu_1_data_master_address_to_slave >> 2;

  //d1_nios_system_clock_8_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_8_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_8_in_end_xfer <= nios_system_clock_8_in_end_xfer;
    end


  //nios_system_clock_8_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_8_in_waits_for_read = nios_system_clock_8_in_in_a_read_cycle & nios_system_clock_8_in_waitrequest_from_sa;

  //nios_system_clock_8_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_8_in_in_a_read_cycle = cpu_1_data_master_granted_nios_system_clock_8_in & cpu_1_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_8_in_in_a_read_cycle;

  //nios_system_clock_8_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_8_in_waits_for_write = nios_system_clock_8_in_in_a_write_cycle & nios_system_clock_8_in_waitrequest_from_sa;

  //nios_system_clock_8_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_8_in_in_a_write_cycle = cpu_1_data_master_granted_nios_system_clock_8_in & cpu_1_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_8_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_8_in_counter = 0;
  //nios_system_clock_8_in_pretend_byte_enable byte enable port mux, which is an e_mux
  assign nios_system_clock_8_in_pretend_byte_enable = (cpu_1_data_master_granted_nios_system_clock_8_in)? cpu_1_data_master_byteenable_nios_system_clock_8_in :
    -1;

  assign {cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_3,
cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_2,
cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_1,
cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_0} = cpu_1_data_master_byteenable;
  assign cpu_1_data_master_byteenable_nios_system_clock_8_in = ((cpu_1_data_master_dbs_address[1 : 0] == 0))? cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_0 :
    ((cpu_1_data_master_dbs_address[1 : 0] == 1))? cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_1 :
    ((cpu_1_data_master_dbs_address[1 : 0] == 2))? cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_2 :
    cpu_1_data_master_byteenable_nios_system_clock_8_in_segment_3;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_8/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_8_out_arbitrator (
                                            // inputs:
                                             clk,
                                             clocks_0_avalon_clocks_slave_readdata_from_sa,
                                             d1_clocks_0_avalon_clocks_slave_end_xfer,
                                             nios_system_clock_8_out_address,
                                             nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave,
                                             nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave,
                                             nios_system_clock_8_out_read,
                                             nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave,
                                             nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave,
                                             nios_system_clock_8_out_write,
                                             nios_system_clock_8_out_writedata,
                                             reset_n,

                                            // outputs:
                                             nios_system_clock_8_out_address_to_slave,
                                             nios_system_clock_8_out_readdata,
                                             nios_system_clock_8_out_reset_n,
                                             nios_system_clock_8_out_waitrequest
                                          )
;

  output           nios_system_clock_8_out_address_to_slave;
  output  [  7: 0] nios_system_clock_8_out_readdata;
  output           nios_system_clock_8_out_reset_n;
  output           nios_system_clock_8_out_waitrequest;
  input            clk;
  input   [  7: 0] clocks_0_avalon_clocks_slave_readdata_from_sa;
  input            d1_clocks_0_avalon_clocks_slave_end_xfer;
  input            nios_system_clock_8_out_address;
  input            nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_8_out_read;
  input            nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_8_out_write;
  input   [  7: 0] nios_system_clock_8_out_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg              nios_system_clock_8_out_address_last_time;
  wire             nios_system_clock_8_out_address_to_slave;
  reg              nios_system_clock_8_out_read_last_time;
  wire    [  7: 0] nios_system_clock_8_out_readdata;
  wire             nios_system_clock_8_out_reset_n;
  wire             nios_system_clock_8_out_run;
  wire             nios_system_clock_8_out_waitrequest;
  reg              nios_system_clock_8_out_write_last_time;
  reg     [  7: 0] nios_system_clock_8_out_writedata_last_time;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave | nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave | ~nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave) & (nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave | ~nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave) & ((~nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave | ~nios_system_clock_8_out_read | (nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave & nios_system_clock_8_out_read))) & ((~nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave | ~(nios_system_clock_8_out_read | nios_system_clock_8_out_write) | (1 & (nios_system_clock_8_out_read | nios_system_clock_8_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_8_out_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_8_out_address_to_slave = nios_system_clock_8_out_address;

  //nios_system_clock_8/out readdata mux, which is an e_mux
  assign nios_system_clock_8_out_readdata = clocks_0_avalon_clocks_slave_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_8_out_waitrequest = ~nios_system_clock_8_out_run;

  //nios_system_clock_8_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_8_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_8_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_8_out_address_last_time <= 0;
      else 
        nios_system_clock_8_out_address_last_time <= nios_system_clock_8_out_address;
    end


  //nios_system_clock_8/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_8_out_waitrequest & (nios_system_clock_8_out_read | nios_system_clock_8_out_write);
    end


  //nios_system_clock_8_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_8_out_address != nios_system_clock_8_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_8_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_8_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_8_out_read_last_time <= 0;
      else 
        nios_system_clock_8_out_read_last_time <= nios_system_clock_8_out_read;
    end


  //nios_system_clock_8_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_8_out_read != nios_system_clock_8_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_8_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_8_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_8_out_write_last_time <= 0;
      else 
        nios_system_clock_8_out_write_last_time <= nios_system_clock_8_out_write;
    end


  //nios_system_clock_8_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_8_out_write != nios_system_clock_8_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_8_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_8_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_8_out_writedata_last_time <= 0;
      else 
        nios_system_clock_8_out_writedata_last_time <= nios_system_clock_8_out_writedata;
    end


  //nios_system_clock_8_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_8_out_writedata != nios_system_clock_8_out_writedata_last_time) & nios_system_clock_8_out_write)
        begin
          $write("%0d ns: nios_system_clock_8_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_9_in_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_0_data_master_address_to_slave,
                                            cpu_0_data_master_byteenable,
                                            cpu_0_data_master_dbs_address,
                                            cpu_0_data_master_dbs_write_8,
                                            cpu_0_data_master_latency_counter,
                                            cpu_0_data_master_read,
                                            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                            cpu_0_data_master_write,
                                            nios_system_clock_9_in_endofpacket,
                                            nios_system_clock_9_in_readdata,
                                            nios_system_clock_9_in_waitrequest,
                                            reset_n,

                                           // outputs:
                                            cpu_0_data_master_byteenable_nios_system_clock_9_in,
                                            cpu_0_data_master_granted_nios_system_clock_9_in,
                                            cpu_0_data_master_qualified_request_nios_system_clock_9_in,
                                            cpu_0_data_master_read_data_valid_nios_system_clock_9_in,
                                            cpu_0_data_master_requests_nios_system_clock_9_in,
                                            d1_nios_system_clock_9_in_end_xfer,
                                            nios_system_clock_9_in_address,
                                            nios_system_clock_9_in_endofpacket_from_sa,
                                            nios_system_clock_9_in_nativeaddress,
                                            nios_system_clock_9_in_read,
                                            nios_system_clock_9_in_readdata_from_sa,
                                            nios_system_clock_9_in_reset_n,
                                            nios_system_clock_9_in_waitrequest_from_sa,
                                            nios_system_clock_9_in_write,
                                            nios_system_clock_9_in_writedata
                                         )
;

  output           cpu_0_data_master_byteenable_nios_system_clock_9_in;
  output           cpu_0_data_master_granted_nios_system_clock_9_in;
  output           cpu_0_data_master_qualified_request_nios_system_clock_9_in;
  output           cpu_0_data_master_read_data_valid_nios_system_clock_9_in;
  output           cpu_0_data_master_requests_nios_system_clock_9_in;
  output           d1_nios_system_clock_9_in_end_xfer;
  output           nios_system_clock_9_in_address;
  output           nios_system_clock_9_in_endofpacket_from_sa;
  output           nios_system_clock_9_in_nativeaddress;
  output           nios_system_clock_9_in_read;
  output  [  7: 0] nios_system_clock_9_in_readdata_from_sa;
  output           nios_system_clock_9_in_reset_n;
  output           nios_system_clock_9_in_waitrequest_from_sa;
  output           nios_system_clock_9_in_write;
  output  [  7: 0] nios_system_clock_9_in_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input   [  1: 0] cpu_0_data_master_dbs_address;
  input   [  7: 0] cpu_0_data_master_dbs_write_8;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input            nios_system_clock_9_in_endofpacket;
  input   [  7: 0] nios_system_clock_9_in_readdata;
  input            nios_system_clock_9_in_waitrequest;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_byteenable_nios_system_clock_9_in;
  wire             cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_0;
  wire             cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_1;
  wire             cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_2;
  wire             cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_3;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_nios_system_clock_9_in;
  wire             cpu_0_data_master_qualified_request_nios_system_clock_9_in;
  wire             cpu_0_data_master_read_data_valid_nios_system_clock_9_in;
  wire             cpu_0_data_master_requests_nios_system_clock_9_in;
  wire             cpu_0_data_master_saved_grant_nios_system_clock_9_in;
  reg              d1_nios_system_clock_9_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_nios_system_clock_9_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             nios_system_clock_9_in_address;
  wire             nios_system_clock_9_in_allgrants;
  wire             nios_system_clock_9_in_allow_new_arb_cycle;
  wire             nios_system_clock_9_in_any_bursting_master_saved_grant;
  wire             nios_system_clock_9_in_any_continuerequest;
  wire             nios_system_clock_9_in_arb_counter_enable;
  reg     [  2: 0] nios_system_clock_9_in_arb_share_counter;
  wire    [  2: 0] nios_system_clock_9_in_arb_share_counter_next_value;
  wire    [  2: 0] nios_system_clock_9_in_arb_share_set_values;
  wire             nios_system_clock_9_in_beginbursttransfer_internal;
  wire             nios_system_clock_9_in_begins_xfer;
  wire             nios_system_clock_9_in_end_xfer;
  wire             nios_system_clock_9_in_endofpacket_from_sa;
  wire             nios_system_clock_9_in_firsttransfer;
  wire             nios_system_clock_9_in_grant_vector;
  wire             nios_system_clock_9_in_in_a_read_cycle;
  wire             nios_system_clock_9_in_in_a_write_cycle;
  wire             nios_system_clock_9_in_master_qreq_vector;
  wire             nios_system_clock_9_in_nativeaddress;
  wire             nios_system_clock_9_in_non_bursting_master_requests;
  wire             nios_system_clock_9_in_pretend_byte_enable;
  wire             nios_system_clock_9_in_read;
  wire    [  7: 0] nios_system_clock_9_in_readdata_from_sa;
  reg              nios_system_clock_9_in_reg_firsttransfer;
  wire             nios_system_clock_9_in_reset_n;
  reg              nios_system_clock_9_in_slavearbiterlockenable;
  wire             nios_system_clock_9_in_slavearbiterlockenable2;
  wire             nios_system_clock_9_in_unreg_firsttransfer;
  wire             nios_system_clock_9_in_waitrequest_from_sa;
  wire             nios_system_clock_9_in_waits_for_read;
  wire             nios_system_clock_9_in_waits_for_write;
  wire             nios_system_clock_9_in_write;
  wire    [  7: 0] nios_system_clock_9_in_writedata;
  wire             wait_for_nios_system_clock_9_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~nios_system_clock_9_in_end_xfer;
    end


  assign nios_system_clock_9_in_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_nios_system_clock_9_in));
  //assign nios_system_clock_9_in_readdata_from_sa = nios_system_clock_9_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_9_in_readdata_from_sa = nios_system_clock_9_in_readdata;

  assign cpu_0_data_master_requests_nios_system_clock_9_in = ({cpu_0_data_master_address_to_slave[24 : 1] , 1'b0} == 25'h19030d8) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //assign nios_system_clock_9_in_waitrequest_from_sa = nios_system_clock_9_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_9_in_waitrequest_from_sa = nios_system_clock_9_in_waitrequest;

  //nios_system_clock_9_in_arb_share_counter set values, which is an e_mux
  assign nios_system_clock_9_in_arb_share_set_values = (cpu_0_data_master_granted_nios_system_clock_9_in)? 4 :
    1;

  //nios_system_clock_9_in_non_bursting_master_requests mux, which is an e_mux
  assign nios_system_clock_9_in_non_bursting_master_requests = cpu_0_data_master_requests_nios_system_clock_9_in;

  //nios_system_clock_9_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign nios_system_clock_9_in_any_bursting_master_saved_grant = 0;

  //nios_system_clock_9_in_arb_share_counter_next_value assignment, which is an e_assign
  assign nios_system_clock_9_in_arb_share_counter_next_value = nios_system_clock_9_in_firsttransfer ? (nios_system_clock_9_in_arb_share_set_values - 1) : |nios_system_clock_9_in_arb_share_counter ? (nios_system_clock_9_in_arb_share_counter - 1) : 0;

  //nios_system_clock_9_in_allgrants all slave grants, which is an e_mux
  assign nios_system_clock_9_in_allgrants = |nios_system_clock_9_in_grant_vector;

  //nios_system_clock_9_in_end_xfer assignment, which is an e_assign
  assign nios_system_clock_9_in_end_xfer = ~(nios_system_clock_9_in_waits_for_read | nios_system_clock_9_in_waits_for_write);

  //end_xfer_arb_share_counter_term_nios_system_clock_9_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_nios_system_clock_9_in = nios_system_clock_9_in_end_xfer & (~nios_system_clock_9_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //nios_system_clock_9_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign nios_system_clock_9_in_arb_counter_enable = (end_xfer_arb_share_counter_term_nios_system_clock_9_in & nios_system_clock_9_in_allgrants) | (end_xfer_arb_share_counter_term_nios_system_clock_9_in & ~nios_system_clock_9_in_non_bursting_master_requests);

  //nios_system_clock_9_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_9_in_arb_share_counter <= 0;
      else if (nios_system_clock_9_in_arb_counter_enable)
          nios_system_clock_9_in_arb_share_counter <= nios_system_clock_9_in_arb_share_counter_next_value;
    end


  //nios_system_clock_9_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_9_in_slavearbiterlockenable <= 0;
      else if ((|nios_system_clock_9_in_master_qreq_vector & end_xfer_arb_share_counter_term_nios_system_clock_9_in) | (end_xfer_arb_share_counter_term_nios_system_clock_9_in & ~nios_system_clock_9_in_non_bursting_master_requests))
          nios_system_clock_9_in_slavearbiterlockenable <= |nios_system_clock_9_in_arb_share_counter_next_value;
    end


  //cpu_0/data_master nios_system_clock_9/in arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = nios_system_clock_9_in_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //nios_system_clock_9_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign nios_system_clock_9_in_slavearbiterlockenable2 = |nios_system_clock_9_in_arb_share_counter_next_value;

  //cpu_0/data_master nios_system_clock_9/in arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = nios_system_clock_9_in_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //nios_system_clock_9_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign nios_system_clock_9_in_any_continuerequest = 1;

  //cpu_0_data_master_continuerequest continued request, which is an e_assign
  assign cpu_0_data_master_continuerequest = 1;

  assign cpu_0_data_master_qualified_request_nios_system_clock_9_in = cpu_0_data_master_requests_nios_system_clock_9_in & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | ((!cpu_0_data_master_byteenable_nios_system_clock_9_in) & cpu_0_data_master_write));
  //local readdatavalid cpu_0_data_master_read_data_valid_nios_system_clock_9_in, which is an e_mux
  assign cpu_0_data_master_read_data_valid_nios_system_clock_9_in = cpu_0_data_master_granted_nios_system_clock_9_in & cpu_0_data_master_read & ~nios_system_clock_9_in_waits_for_read;

  //nios_system_clock_9_in_writedata mux, which is an e_mux
  assign nios_system_clock_9_in_writedata = cpu_0_data_master_dbs_write_8;

  //assign nios_system_clock_9_in_endofpacket_from_sa = nios_system_clock_9_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign nios_system_clock_9_in_endofpacket_from_sa = nios_system_clock_9_in_endofpacket;

  //master is always granted when requested
  assign cpu_0_data_master_granted_nios_system_clock_9_in = cpu_0_data_master_qualified_request_nios_system_clock_9_in;

  //cpu_0/data_master saved-grant nios_system_clock_9/in, which is an e_assign
  assign cpu_0_data_master_saved_grant_nios_system_clock_9_in = cpu_0_data_master_requests_nios_system_clock_9_in;

  //allow new arb cycle for nios_system_clock_9/in, which is an e_assign
  assign nios_system_clock_9_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign nios_system_clock_9_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign nios_system_clock_9_in_master_qreq_vector = 1;

  //nios_system_clock_9_in_reset_n assignment, which is an e_assign
  assign nios_system_clock_9_in_reset_n = reset_n;

  //nios_system_clock_9_in_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_9_in_firsttransfer = nios_system_clock_9_in_begins_xfer ? nios_system_clock_9_in_unreg_firsttransfer : nios_system_clock_9_in_reg_firsttransfer;

  //nios_system_clock_9_in_unreg_firsttransfer first transaction, which is an e_assign
  assign nios_system_clock_9_in_unreg_firsttransfer = ~(nios_system_clock_9_in_slavearbiterlockenable & nios_system_clock_9_in_any_continuerequest);

  //nios_system_clock_9_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_9_in_reg_firsttransfer <= 1'b1;
      else if (nios_system_clock_9_in_begins_xfer)
          nios_system_clock_9_in_reg_firsttransfer <= nios_system_clock_9_in_unreg_firsttransfer;
    end


  //nios_system_clock_9_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign nios_system_clock_9_in_beginbursttransfer_internal = nios_system_clock_9_in_begins_xfer;

  //nios_system_clock_9_in_read assignment, which is an e_mux
  assign nios_system_clock_9_in_read = cpu_0_data_master_granted_nios_system_clock_9_in & cpu_0_data_master_read;

  //nios_system_clock_9_in_write assignment, which is an e_mux
  assign nios_system_clock_9_in_write = ((cpu_0_data_master_granted_nios_system_clock_9_in & cpu_0_data_master_write)) & nios_system_clock_9_in_pretend_byte_enable;

  //nios_system_clock_9_in_address mux, which is an e_mux
  assign nios_system_clock_9_in_address = {cpu_0_data_master_address_to_slave >> 2,
    cpu_0_data_master_dbs_address[1 : 0]};

  //slaveid nios_system_clock_9_in_nativeaddress nativeaddress mux, which is an e_mux
  assign nios_system_clock_9_in_nativeaddress = cpu_0_data_master_address_to_slave >> 2;

  //d1_nios_system_clock_9_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_nios_system_clock_9_in_end_xfer <= 1;
      else 
        d1_nios_system_clock_9_in_end_xfer <= nios_system_clock_9_in_end_xfer;
    end


  //nios_system_clock_9_in_waits_for_read in a cycle, which is an e_mux
  assign nios_system_clock_9_in_waits_for_read = nios_system_clock_9_in_in_a_read_cycle & nios_system_clock_9_in_waitrequest_from_sa;

  //nios_system_clock_9_in_in_a_read_cycle assignment, which is an e_assign
  assign nios_system_clock_9_in_in_a_read_cycle = cpu_0_data_master_granted_nios_system_clock_9_in & cpu_0_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = nios_system_clock_9_in_in_a_read_cycle;

  //nios_system_clock_9_in_waits_for_write in a cycle, which is an e_mux
  assign nios_system_clock_9_in_waits_for_write = nios_system_clock_9_in_in_a_write_cycle & nios_system_clock_9_in_waitrequest_from_sa;

  //nios_system_clock_9_in_in_a_write_cycle assignment, which is an e_assign
  assign nios_system_clock_9_in_in_a_write_cycle = cpu_0_data_master_granted_nios_system_clock_9_in & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = nios_system_clock_9_in_in_a_write_cycle;

  assign wait_for_nios_system_clock_9_in_counter = 0;
  //nios_system_clock_9_in_pretend_byte_enable byte enable port mux, which is an e_mux
  assign nios_system_clock_9_in_pretend_byte_enable = (cpu_0_data_master_granted_nios_system_clock_9_in)? cpu_0_data_master_byteenable_nios_system_clock_9_in :
    -1;

  assign {cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_3,
cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_2,
cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_1,
cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_0} = cpu_0_data_master_byteenable;
  assign cpu_0_data_master_byteenable_nios_system_clock_9_in = ((cpu_0_data_master_dbs_address[1 : 0] == 0))? cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_0 :
    ((cpu_0_data_master_dbs_address[1 : 0] == 1))? cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_1 :
    ((cpu_0_data_master_dbs_address[1 : 0] == 2))? cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_2 :
    cpu_0_data_master_byteenable_nios_system_clock_9_in_segment_3;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_9/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_clock_9_out_arbitrator (
                                            // inputs:
                                             clk,
                                             clocks_0_avalon_clocks_slave_readdata_from_sa,
                                             d1_clocks_0_avalon_clocks_slave_end_xfer,
                                             nios_system_clock_9_out_address,
                                             nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave,
                                             nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave,
                                             nios_system_clock_9_out_read,
                                             nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave,
                                             nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave,
                                             nios_system_clock_9_out_write,
                                             nios_system_clock_9_out_writedata,
                                             reset_n,

                                            // outputs:
                                             nios_system_clock_9_out_address_to_slave,
                                             nios_system_clock_9_out_readdata,
                                             nios_system_clock_9_out_reset_n,
                                             nios_system_clock_9_out_waitrequest
                                          )
;

  output           nios_system_clock_9_out_address_to_slave;
  output  [  7: 0] nios_system_clock_9_out_readdata;
  output           nios_system_clock_9_out_reset_n;
  output           nios_system_clock_9_out_waitrequest;
  input            clk;
  input   [  7: 0] clocks_0_avalon_clocks_slave_readdata_from_sa;
  input            d1_clocks_0_avalon_clocks_slave_end_xfer;
  input            nios_system_clock_9_out_address;
  input            nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_9_out_read;
  input            nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave;
  input            nios_system_clock_9_out_write;
  input   [  7: 0] nios_system_clock_9_out_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg              nios_system_clock_9_out_address_last_time;
  wire             nios_system_clock_9_out_address_to_slave;
  reg              nios_system_clock_9_out_read_last_time;
  wire    [  7: 0] nios_system_clock_9_out_readdata;
  wire             nios_system_clock_9_out_reset_n;
  wire             nios_system_clock_9_out_run;
  wire             nios_system_clock_9_out_waitrequest;
  reg              nios_system_clock_9_out_write_last_time;
  reg     [  7: 0] nios_system_clock_9_out_writedata_last_time;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave | nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave | ~nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave) & (nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave | ~nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave) & ((~nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave | ~nios_system_clock_9_out_read | (nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave & nios_system_clock_9_out_read))) & ((~nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave | ~(nios_system_clock_9_out_read | nios_system_clock_9_out_write) | (1 & (nios_system_clock_9_out_read | nios_system_clock_9_out_write))));

  //cascaded wait assignment, which is an e_assign
  assign nios_system_clock_9_out_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign nios_system_clock_9_out_address_to_slave = nios_system_clock_9_out_address;

  //nios_system_clock_9/out readdata mux, which is an e_mux
  assign nios_system_clock_9_out_readdata = clocks_0_avalon_clocks_slave_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign nios_system_clock_9_out_waitrequest = ~nios_system_clock_9_out_run;

  //nios_system_clock_9_out_reset_n assignment, which is an e_assign
  assign nios_system_clock_9_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //nios_system_clock_9_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_9_out_address_last_time <= 0;
      else 
        nios_system_clock_9_out_address_last_time <= nios_system_clock_9_out_address;
    end


  //nios_system_clock_9/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= nios_system_clock_9_out_waitrequest & (nios_system_clock_9_out_read | nios_system_clock_9_out_write);
    end


  //nios_system_clock_9_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_9_out_address != nios_system_clock_9_out_address_last_time))
        begin
          $write("%0d ns: nios_system_clock_9_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_9_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_9_out_read_last_time <= 0;
      else 
        nios_system_clock_9_out_read_last_time <= nios_system_clock_9_out_read;
    end


  //nios_system_clock_9_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_9_out_read != nios_system_clock_9_out_read_last_time))
        begin
          $write("%0d ns: nios_system_clock_9_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_9_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_9_out_write_last_time <= 0;
      else 
        nios_system_clock_9_out_write_last_time <= nios_system_clock_9_out_write;
    end


  //nios_system_clock_9_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_9_out_write != nios_system_clock_9_out_write_last_time))
        begin
          $write("%0d ns: nios_system_clock_9_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //nios_system_clock_9_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          nios_system_clock_9_out_writedata_last_time <= 0;
      else 
        nios_system_clock_9_out_writedata_last_time <= nios_system_clock_9_out_writedata;
    end


  //nios_system_clock_9_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (nios_system_clock_9_out_writedata != nios_system_clock_9_out_writedata_last_time) & nios_system_clock_9_out_write)
        begin
          $write("%0d ns: nios_system_clock_9_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module onchip_memory2_0_s1_arbitrator (
                                        // inputs:
                                         clk,
                                         cpu_0_data_master_address_to_slave,
                                         cpu_0_data_master_byteenable,
                                         cpu_0_data_master_latency_counter,
                                         cpu_0_data_master_read,
                                         cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_0_data_master_write,
                                         cpu_0_data_master_writedata,
                                         cpu_0_instruction_master_address_to_slave,
                                         cpu_0_instruction_master_latency_counter,
                                         cpu_0_instruction_master_read,
                                         cpu_1_data_master_address_to_slave,
                                         cpu_1_data_master_byteenable,
                                         cpu_1_data_master_latency_counter,
                                         cpu_1_data_master_read,
                                         cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_1_data_master_write,
                                         cpu_1_data_master_writedata,
                                         cpu_1_instruction_master_address_to_slave,
                                         cpu_1_instruction_master_latency_counter,
                                         cpu_1_instruction_master_read,
                                         cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_2_data_master_address_to_slave,
                                         cpu_2_data_master_byteenable,
                                         cpu_2_data_master_latency_counter,
                                         cpu_2_data_master_read,
                                         cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_2_data_master_write,
                                         cpu_2_data_master_writedata,
                                         cpu_2_instruction_master_address_to_slave,
                                         cpu_2_instruction_master_latency_counter,
                                         cpu_2_instruction_master_read,
                                         cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_3_data_master_address_to_slave,
                                         cpu_3_data_master_byteenable,
                                         cpu_3_data_master_latency_counter,
                                         cpu_3_data_master_read,
                                         cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_3_data_master_write,
                                         cpu_3_data_master_writedata,
                                         cpu_3_instruction_master_address_to_slave,
                                         cpu_3_instruction_master_latency_counter,
                                         cpu_3_instruction_master_read,
                                         cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         onchip_memory2_0_s1_readdata,
                                         reset_n,

                                        // outputs:
                                         cpu_0_data_master_granted_onchip_memory2_0_s1,
                                         cpu_0_data_master_qualified_request_onchip_memory2_0_s1,
                                         cpu_0_data_master_read_data_valid_onchip_memory2_0_s1,
                                         cpu_0_data_master_requests_onchip_memory2_0_s1,
                                         cpu_0_instruction_master_granted_onchip_memory2_0_s1,
                                         cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1,
                                         cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1,
                                         cpu_0_instruction_master_requests_onchip_memory2_0_s1,
                                         cpu_1_data_master_granted_onchip_memory2_0_s1,
                                         cpu_1_data_master_qualified_request_onchip_memory2_0_s1,
                                         cpu_1_data_master_read_data_valid_onchip_memory2_0_s1,
                                         cpu_1_data_master_requests_onchip_memory2_0_s1,
                                         cpu_1_instruction_master_granted_onchip_memory2_0_s1,
                                         cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1,
                                         cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1,
                                         cpu_1_instruction_master_requests_onchip_memory2_0_s1,
                                         cpu_2_data_master_granted_onchip_memory2_0_s1,
                                         cpu_2_data_master_qualified_request_onchip_memory2_0_s1,
                                         cpu_2_data_master_read_data_valid_onchip_memory2_0_s1,
                                         cpu_2_data_master_requests_onchip_memory2_0_s1,
                                         cpu_2_instruction_master_granted_onchip_memory2_0_s1,
                                         cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1,
                                         cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1,
                                         cpu_2_instruction_master_requests_onchip_memory2_0_s1,
                                         cpu_3_data_master_granted_onchip_memory2_0_s1,
                                         cpu_3_data_master_qualified_request_onchip_memory2_0_s1,
                                         cpu_3_data_master_read_data_valid_onchip_memory2_0_s1,
                                         cpu_3_data_master_requests_onchip_memory2_0_s1,
                                         cpu_3_instruction_master_granted_onchip_memory2_0_s1,
                                         cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1,
                                         cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1,
                                         cpu_3_instruction_master_requests_onchip_memory2_0_s1,
                                         d1_onchip_memory2_0_s1_end_xfer,
                                         onchip_memory2_0_s1_address,
                                         onchip_memory2_0_s1_byteenable,
                                         onchip_memory2_0_s1_chipselect,
                                         onchip_memory2_0_s1_clken,
                                         onchip_memory2_0_s1_readdata_from_sa,
                                         onchip_memory2_0_s1_reset,
                                         onchip_memory2_0_s1_write,
                                         onchip_memory2_0_s1_writedata
                                      )
;

  output           cpu_0_data_master_granted_onchip_memory2_0_s1;
  output           cpu_0_data_master_qualified_request_onchip_memory2_0_s1;
  output           cpu_0_data_master_read_data_valid_onchip_memory2_0_s1;
  output           cpu_0_data_master_requests_onchip_memory2_0_s1;
  output           cpu_0_instruction_master_granted_onchip_memory2_0_s1;
  output           cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1;
  output           cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1;
  output           cpu_0_instruction_master_requests_onchip_memory2_0_s1;
  output           cpu_1_data_master_granted_onchip_memory2_0_s1;
  output           cpu_1_data_master_qualified_request_onchip_memory2_0_s1;
  output           cpu_1_data_master_read_data_valid_onchip_memory2_0_s1;
  output           cpu_1_data_master_requests_onchip_memory2_0_s1;
  output           cpu_1_instruction_master_granted_onchip_memory2_0_s1;
  output           cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1;
  output           cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1;
  output           cpu_1_instruction_master_requests_onchip_memory2_0_s1;
  output           cpu_2_data_master_granted_onchip_memory2_0_s1;
  output           cpu_2_data_master_qualified_request_onchip_memory2_0_s1;
  output           cpu_2_data_master_read_data_valid_onchip_memory2_0_s1;
  output           cpu_2_data_master_requests_onchip_memory2_0_s1;
  output           cpu_2_instruction_master_granted_onchip_memory2_0_s1;
  output           cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1;
  output           cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1;
  output           cpu_2_instruction_master_requests_onchip_memory2_0_s1;
  output           cpu_3_data_master_granted_onchip_memory2_0_s1;
  output           cpu_3_data_master_qualified_request_onchip_memory2_0_s1;
  output           cpu_3_data_master_read_data_valid_onchip_memory2_0_s1;
  output           cpu_3_data_master_requests_onchip_memory2_0_s1;
  output           cpu_3_instruction_master_granted_onchip_memory2_0_s1;
  output           cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1;
  output           cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1;
  output           cpu_3_instruction_master_requests_onchip_memory2_0_s1;
  output           d1_onchip_memory2_0_s1_end_xfer;
  output  [  6: 0] onchip_memory2_0_s1_address;
  output  [  3: 0] onchip_memory2_0_s1_byteenable;
  output           onchip_memory2_0_s1_chipselect;
  output           onchip_memory2_0_s1_clken;
  output  [ 31: 0] onchip_memory2_0_s1_readdata_from_sa;
  output           onchip_memory2_0_s1_reset;
  output           onchip_memory2_0_s1_write;
  output  [ 31: 0] onchip_memory2_0_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input            cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input   [  3: 0] cpu_1_data_master_byteenable;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_1_instruction_master_address_to_slave;
  input            cpu_1_instruction_master_latency_counter;
  input            cpu_1_instruction_master_read;
  input            cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input   [  3: 0] cpu_2_data_master_byteenable;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_2_instruction_master_address_to_slave;
  input            cpu_2_instruction_master_latency_counter;
  input            cpu_2_instruction_master_read;
  input            cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input   [  3: 0] cpu_3_data_master_byteenable;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 24: 0] cpu_3_instruction_master_address_to_slave;
  input            cpu_3_instruction_master_latency_counter;
  input            cpu_3_instruction_master_read;
  input            cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 31: 0] onchip_memory2_0_s1_readdata;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_onchip_memory2_0_s1;
  wire             cpu_0_data_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_0_s1;
  reg              cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in;
  wire             cpu_0_data_master_requests_onchip_memory2_0_s1;
  wire             cpu_0_data_master_saved_grant_onchip_memory2_0_s1;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_onchip_memory2_0_s1;
  wire             cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1;
  reg              cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in;
  wire             cpu_0_instruction_master_requests_onchip_memory2_0_s1;
  wire             cpu_0_instruction_master_saved_grant_onchip_memory2_0_s1;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_onchip_memory2_0_s1;
  wire             cpu_1_data_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_0_s1;
  reg              cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in;
  wire             cpu_1_data_master_requests_onchip_memory2_0_s1;
  wire             cpu_1_data_master_saved_grant_onchip_memory2_0_s1;
  wire             cpu_1_instruction_master_arbiterlock;
  wire             cpu_1_instruction_master_arbiterlock2;
  wire             cpu_1_instruction_master_continuerequest;
  wire             cpu_1_instruction_master_granted_onchip_memory2_0_s1;
  wire             cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1;
  reg              cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in;
  wire             cpu_1_instruction_master_requests_onchip_memory2_0_s1;
  wire             cpu_1_instruction_master_saved_grant_onchip_memory2_0_s1;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_onchip_memory2_0_s1;
  wire             cpu_2_data_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_0_s1;
  reg              cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in;
  wire             cpu_2_data_master_requests_onchip_memory2_0_s1;
  wire             cpu_2_data_master_saved_grant_onchip_memory2_0_s1;
  wire             cpu_2_instruction_master_arbiterlock;
  wire             cpu_2_instruction_master_arbiterlock2;
  wire             cpu_2_instruction_master_continuerequest;
  wire             cpu_2_instruction_master_granted_onchip_memory2_0_s1;
  wire             cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1;
  reg              cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in;
  wire             cpu_2_instruction_master_requests_onchip_memory2_0_s1;
  wire             cpu_2_instruction_master_saved_grant_onchip_memory2_0_s1;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_onchip_memory2_0_s1;
  wire             cpu_3_data_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_0_s1;
  reg              cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in;
  wire             cpu_3_data_master_requests_onchip_memory2_0_s1;
  wire             cpu_3_data_master_saved_grant_onchip_memory2_0_s1;
  wire             cpu_3_instruction_master_arbiterlock;
  wire             cpu_3_instruction_master_arbiterlock2;
  wire             cpu_3_instruction_master_continuerequest;
  wire             cpu_3_instruction_master_granted_onchip_memory2_0_s1;
  wire             cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1;
  reg              cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in;
  wire             cpu_3_instruction_master_requests_onchip_memory2_0_s1;
  wire             cpu_3_instruction_master_saved_grant_onchip_memory2_0_s1;
  reg              d1_onchip_memory2_0_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_onchip_memory2_0_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_0_s1;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_0_s1;
  reg              last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_0_s1;
  reg              last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_0_s1;
  reg              last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_0_s1;
  reg              last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_0_s1;
  reg              last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_0_s1;
  reg              last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_0_s1;
  wire    [  6: 0] onchip_memory2_0_s1_address;
  wire             onchip_memory2_0_s1_allgrants;
  wire             onchip_memory2_0_s1_allow_new_arb_cycle;
  wire             onchip_memory2_0_s1_any_bursting_master_saved_grant;
  wire             onchip_memory2_0_s1_any_continuerequest;
  reg     [  7: 0] onchip_memory2_0_s1_arb_addend;
  wire             onchip_memory2_0_s1_arb_counter_enable;
  reg     [  2: 0] onchip_memory2_0_s1_arb_share_counter;
  wire    [  2: 0] onchip_memory2_0_s1_arb_share_counter_next_value;
  wire    [  2: 0] onchip_memory2_0_s1_arb_share_set_values;
  wire    [  7: 0] onchip_memory2_0_s1_arb_winner;
  wire             onchip_memory2_0_s1_arbitration_holdoff_internal;
  wire             onchip_memory2_0_s1_beginbursttransfer_internal;
  wire             onchip_memory2_0_s1_begins_xfer;
  wire    [  3: 0] onchip_memory2_0_s1_byteenable;
  wire             onchip_memory2_0_s1_chipselect;
  wire    [ 15: 0] onchip_memory2_0_s1_chosen_master_double_vector;
  wire    [  7: 0] onchip_memory2_0_s1_chosen_master_rot_left;
  wire             onchip_memory2_0_s1_clken;
  wire             onchip_memory2_0_s1_end_xfer;
  wire             onchip_memory2_0_s1_firsttransfer;
  wire    [  7: 0] onchip_memory2_0_s1_grant_vector;
  wire             onchip_memory2_0_s1_in_a_read_cycle;
  wire             onchip_memory2_0_s1_in_a_write_cycle;
  wire    [  7: 0] onchip_memory2_0_s1_master_qreq_vector;
  wire             onchip_memory2_0_s1_non_bursting_master_requests;
  wire    [ 31: 0] onchip_memory2_0_s1_readdata_from_sa;
  reg              onchip_memory2_0_s1_reg_firsttransfer;
  wire             onchip_memory2_0_s1_reset;
  reg     [  7: 0] onchip_memory2_0_s1_saved_chosen_master_vector;
  reg              onchip_memory2_0_s1_slavearbiterlockenable;
  wire             onchip_memory2_0_s1_slavearbiterlockenable2;
  wire             onchip_memory2_0_s1_unreg_firsttransfer;
  wire             onchip_memory2_0_s1_waits_for_read;
  wire             onchip_memory2_0_s1_waits_for_write;
  wire             onchip_memory2_0_s1_write;
  wire    [ 31: 0] onchip_memory2_0_s1_writedata;
  wire             p1_cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             p1_cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             p1_cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             p1_cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire             p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_0_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_0_s1_from_cpu_0_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_0_s1_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_0_s1_from_cpu_1_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_0_s1_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_0_s1_from_cpu_2_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_0_s1_from_cpu_3_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_0_s1_from_cpu_3_instruction_master;
  wire             wait_for_onchip_memory2_0_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~onchip_memory2_0_s1_end_xfer;
    end


  assign onchip_memory2_0_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_onchip_memory2_0_s1 | cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1 | cpu_1_data_master_qualified_request_onchip_memory2_0_s1 | cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1 | cpu_2_data_master_qualified_request_onchip_memory2_0_s1 | cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1 | cpu_3_data_master_qualified_request_onchip_memory2_0_s1 | cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1));
  //assign onchip_memory2_0_s1_readdata_from_sa = onchip_memory2_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign onchip_memory2_0_s1_readdata_from_sa = onchip_memory2_0_s1_readdata;

  assign cpu_0_data_master_requests_onchip_memory2_0_s1 = ({cpu_0_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h3000) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //onchip_memory2_0_s1_arb_share_counter set values, which is an e_mux
  assign onchip_memory2_0_s1_arb_share_set_values = 1;

  //onchip_memory2_0_s1_non_bursting_master_requests mux, which is an e_mux
  assign onchip_memory2_0_s1_non_bursting_master_requests = cpu_0_data_master_requests_onchip_memory2_0_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_1_data_master_requests_onchip_memory2_0_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_2_data_master_requests_onchip_memory2_0_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_3_data_master_requests_onchip_memory2_0_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_0_data_master_requests_onchip_memory2_0_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_1_data_master_requests_onchip_memory2_0_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_2_data_master_requests_onchip_memory2_0_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_3_data_master_requests_onchip_memory2_0_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_0_data_master_requests_onchip_memory2_0_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_1_data_master_requests_onchip_memory2_0_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_2_data_master_requests_onchip_memory2_0_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_3_data_master_requests_onchip_memory2_0_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_0_data_master_requests_onchip_memory2_0_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_1_data_master_requests_onchip_memory2_0_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_2_data_master_requests_onchip_memory2_0_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_3_data_master_requests_onchip_memory2_0_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_0_data_master_requests_onchip_memory2_0_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_1_data_master_requests_onchip_memory2_0_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_2_data_master_requests_onchip_memory2_0_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_3_data_master_requests_onchip_memory2_0_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_0_data_master_requests_onchip_memory2_0_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_1_data_master_requests_onchip_memory2_0_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_2_data_master_requests_onchip_memory2_0_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_3_data_master_requests_onchip_memory2_0_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_0_data_master_requests_onchip_memory2_0_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_1_data_master_requests_onchip_memory2_0_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_2_data_master_requests_onchip_memory2_0_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_3_data_master_requests_onchip_memory2_0_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_0_data_master_requests_onchip_memory2_0_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_1_data_master_requests_onchip_memory2_0_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_2_data_master_requests_onchip_memory2_0_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_0_s1 |
    cpu_3_data_master_requests_onchip_memory2_0_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_0_s1;

  //onchip_memory2_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign onchip_memory2_0_s1_any_bursting_master_saved_grant = 0;

  //onchip_memory2_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign onchip_memory2_0_s1_arb_share_counter_next_value = onchip_memory2_0_s1_firsttransfer ? (onchip_memory2_0_s1_arb_share_set_values - 1) : |onchip_memory2_0_s1_arb_share_counter ? (onchip_memory2_0_s1_arb_share_counter - 1) : 0;

  //onchip_memory2_0_s1_allgrants all slave grants, which is an e_mux
  assign onchip_memory2_0_s1_allgrants = (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector) |
    (|onchip_memory2_0_s1_grant_vector);

  //onchip_memory2_0_s1_end_xfer assignment, which is an e_assign
  assign onchip_memory2_0_s1_end_xfer = ~(onchip_memory2_0_s1_waits_for_read | onchip_memory2_0_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_onchip_memory2_0_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_onchip_memory2_0_s1 = onchip_memory2_0_s1_end_xfer & (~onchip_memory2_0_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //onchip_memory2_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign onchip_memory2_0_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_onchip_memory2_0_s1 & onchip_memory2_0_s1_allgrants) | (end_xfer_arb_share_counter_term_onchip_memory2_0_s1 & ~onchip_memory2_0_s1_non_bursting_master_requests);

  //onchip_memory2_0_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_0_s1_arb_share_counter <= 0;
      else if (onchip_memory2_0_s1_arb_counter_enable)
          onchip_memory2_0_s1_arb_share_counter <= onchip_memory2_0_s1_arb_share_counter_next_value;
    end


  //onchip_memory2_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_0_s1_slavearbiterlockenable <= 0;
      else if ((|onchip_memory2_0_s1_master_qreq_vector & end_xfer_arb_share_counter_term_onchip_memory2_0_s1) | (end_xfer_arb_share_counter_term_onchip_memory2_0_s1 & ~onchip_memory2_0_s1_non_bursting_master_requests))
          onchip_memory2_0_s1_slavearbiterlockenable <= |onchip_memory2_0_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master onchip_memory2_0/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = onchip_memory2_0_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //onchip_memory2_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign onchip_memory2_0_s1_slavearbiterlockenable2 = |onchip_memory2_0_s1_arb_share_counter_next_value;

  //cpu_0/data_master onchip_memory2_0/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = onchip_memory2_0_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master onchip_memory2_0/s1 arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = onchip_memory2_0_s1_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master onchip_memory2_0/s1 arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = onchip_memory2_0_s1_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted onchip_memory2_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_0_s1 <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_0_s1 <= cpu_0_instruction_master_saved_grant_onchip_memory2_0_s1 ? 1 : (onchip_memory2_0_s1_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_onchip_memory2_0_s1) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_0_s1;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_0_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_0_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_0_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_0_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_0_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_0_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_0_instruction_master_requests_onchip_memory2_0_s1);

  //onchip_memory2_0_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign onchip_memory2_0_s1_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest;

  //cpu_1/data_master onchip_memory2_0/s1 arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = onchip_memory2_0_s1_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master onchip_memory2_0/s1 arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = onchip_memory2_0_s1_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted onchip_memory2_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_0_s1 <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_0_s1 <= cpu_1_data_master_saved_grant_onchip_memory2_0_s1 ? 1 : (onchip_memory2_0_s1_arbitration_holdoff_internal | ~cpu_1_data_master_requests_onchip_memory2_0_s1) ? 0 : last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_0_s1;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_0_s1 & cpu_1_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_0_s1 & cpu_1_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_0_s1 & cpu_1_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_0_s1 & cpu_1_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_0_s1 & cpu_1_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_0_s1 & cpu_1_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_0_s1 & cpu_1_data_master_requests_onchip_memory2_0_s1);

  //cpu_1/instruction_master onchip_memory2_0/s1 arbiterlock, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock = onchip_memory2_0_s1_slavearbiterlockenable & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master onchip_memory2_0/s1 arbiterlock2, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock2 = onchip_memory2_0_s1_slavearbiterlockenable2 & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master granted onchip_memory2_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_0_s1 <= 0;
      else 
        last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_0_s1 <= cpu_1_instruction_master_saved_grant_onchip_memory2_0_s1 ? 1 : (onchip_memory2_0_s1_arbitration_holdoff_internal | ~cpu_1_instruction_master_requests_onchip_memory2_0_s1) ? 0 : last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_0_s1;
    end


  //cpu_1_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_1_instruction_master_continuerequest = (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_1_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_1_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_1_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_1_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_1_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_1_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_1_instruction_master_requests_onchip_memory2_0_s1);

  //cpu_2/data_master onchip_memory2_0/s1 arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = onchip_memory2_0_s1_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master onchip_memory2_0/s1 arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = onchip_memory2_0_s1_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted onchip_memory2_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_0_s1 <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_0_s1 <= cpu_2_data_master_saved_grant_onchip_memory2_0_s1 ? 1 : (onchip_memory2_0_s1_arbitration_holdoff_internal | ~cpu_2_data_master_requests_onchip_memory2_0_s1) ? 0 : last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_0_s1;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_0_s1 & cpu_2_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_0_s1 & cpu_2_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_0_s1 & cpu_2_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_0_s1 & cpu_2_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_0_s1 & cpu_2_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_0_s1 & cpu_2_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_0_s1 & cpu_2_data_master_requests_onchip_memory2_0_s1);

  //cpu_2/instruction_master onchip_memory2_0/s1 arbiterlock, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock = onchip_memory2_0_s1_slavearbiterlockenable & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master onchip_memory2_0/s1 arbiterlock2, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock2 = onchip_memory2_0_s1_slavearbiterlockenable2 & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master granted onchip_memory2_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_0_s1 <= 0;
      else 
        last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_0_s1 <= cpu_2_instruction_master_saved_grant_onchip_memory2_0_s1 ? 1 : (onchip_memory2_0_s1_arbitration_holdoff_internal | ~cpu_2_instruction_master_requests_onchip_memory2_0_s1) ? 0 : last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_0_s1;
    end


  //cpu_2_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_2_instruction_master_continuerequest = (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_2_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_2_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_2_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_2_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_2_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_2_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_2_instruction_master_requests_onchip_memory2_0_s1);

  //cpu_3/data_master onchip_memory2_0/s1 arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = onchip_memory2_0_s1_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master onchip_memory2_0/s1 arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = onchip_memory2_0_s1_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted onchip_memory2_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_0_s1 <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_0_s1 <= cpu_3_data_master_saved_grant_onchip_memory2_0_s1 ? 1 : (onchip_memory2_0_s1_arbitration_holdoff_internal | ~cpu_3_data_master_requests_onchip_memory2_0_s1) ? 0 : last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_0_s1;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_0_s1 & cpu_3_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_0_s1 & cpu_3_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_0_s1 & cpu_3_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_0_s1 & cpu_3_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_0_s1 & cpu_3_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_0_s1 & cpu_3_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_0_s1 & cpu_3_data_master_requests_onchip_memory2_0_s1);

  //cpu_3/instruction_master onchip_memory2_0/s1 arbiterlock, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock = onchip_memory2_0_s1_slavearbiterlockenable & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master onchip_memory2_0/s1 arbiterlock2, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock2 = onchip_memory2_0_s1_slavearbiterlockenable2 & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master granted onchip_memory2_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_0_s1 <= 0;
      else 
        last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_0_s1 <= cpu_3_instruction_master_saved_grant_onchip_memory2_0_s1 ? 1 : (onchip_memory2_0_s1_arbitration_holdoff_internal | ~cpu_3_instruction_master_requests_onchip_memory2_0_s1) ? 0 : last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_0_s1;
    end


  //cpu_3_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_3_instruction_master_continuerequest = (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_3_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_3_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_3_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_3_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_3_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_3_instruction_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_0_s1 & cpu_3_instruction_master_requests_onchip_memory2_0_s1);

  assign cpu_0_data_master_qualified_request_onchip_memory2_0_s1 = cpu_0_data_master_requests_onchip_memory2_0_s1 & ~((cpu_0_data_master_read & ((1 < cpu_0_data_master_latency_counter) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in = cpu_0_data_master_granted_onchip_memory2_0_s1 & cpu_0_data_master_read & ~onchip_memory2_0_s1_waits_for_read;

  //shift register p1 cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register = {cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register, cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in};

  //cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register <= 0;
      else 
        cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register <= p1_cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
    end


  //local readdatavalid cpu_0_data_master_read_data_valid_onchip_memory2_0_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_onchip_memory2_0_s1 = cpu_0_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;

  //onchip_memory2_0_s1_writedata mux, which is an e_mux
  assign onchip_memory2_0_s1_writedata = (cpu_0_data_master_granted_onchip_memory2_0_s1)? cpu_0_data_master_writedata :
    (cpu_1_data_master_granted_onchip_memory2_0_s1)? cpu_1_data_master_writedata :
    (cpu_2_data_master_granted_onchip_memory2_0_s1)? cpu_2_data_master_writedata :
    cpu_3_data_master_writedata;

  //mux onchip_memory2_0_s1_clken, which is an e_mux
  assign onchip_memory2_0_s1_clken = 1'b1;

  assign cpu_0_instruction_master_requests_onchip_memory2_0_s1 = (({cpu_0_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h3000) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted onchip_memory2_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_0_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_0_s1 <= cpu_0_data_master_saved_grant_onchip_memory2_0_s1 ? 1 : (onchip_memory2_0_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_onchip_memory2_0_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_0_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_0_s1 & cpu_0_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_0_s1 & cpu_0_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_0_s1 & cpu_0_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_0_s1 & cpu_0_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_0_s1 & cpu_0_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_0_s1 & cpu_0_data_master_requests_onchip_memory2_0_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_0_s1 & cpu_0_data_master_requests_onchip_memory2_0_s1);

  assign cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1 = cpu_0_instruction_master_requests_onchip_memory2_0_s1 & ~((cpu_0_instruction_master_read & ((1 < cpu_0_instruction_master_latency_counter))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in = cpu_0_instruction_master_granted_onchip_memory2_0_s1 & cpu_0_instruction_master_read & ~onchip_memory2_0_s1_waits_for_read;

  //shift register p1 cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register = {cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register, cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in};

  //cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register <= 0;
      else 
        cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register <= p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
    end


  //local readdatavalid cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1 = cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;

  assign cpu_1_data_master_requests_onchip_memory2_0_s1 = ({cpu_1_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h3000) & (cpu_1_data_master_read | cpu_1_data_master_write);
  assign cpu_1_data_master_qualified_request_onchip_memory2_0_s1 = cpu_1_data_master_requests_onchip_memory2_0_s1 & ~((cpu_1_data_master_read & ((1 < cpu_1_data_master_latency_counter) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in = cpu_1_data_master_granted_onchip_memory2_0_s1 & cpu_1_data_master_read & ~onchip_memory2_0_s1_waits_for_read;

  //shift register p1 cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register = {cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register, cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in};

  //cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register <= 0;
      else 
        cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register <= p1_cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
    end


  //local readdatavalid cpu_1_data_master_read_data_valid_onchip_memory2_0_s1, which is an e_mux
  assign cpu_1_data_master_read_data_valid_onchip_memory2_0_s1 = cpu_1_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;

  assign cpu_1_instruction_master_requests_onchip_memory2_0_s1 = (({cpu_1_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h3000) & (cpu_1_instruction_master_read)) & cpu_1_instruction_master_read;
  assign cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1 = cpu_1_instruction_master_requests_onchip_memory2_0_s1 & ~((cpu_1_instruction_master_read & ((1 < cpu_1_instruction_master_latency_counter) | (|cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in = cpu_1_instruction_master_granted_onchip_memory2_0_s1 & cpu_1_instruction_master_read & ~onchip_memory2_0_s1_waits_for_read;

  //shift register p1 cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register = {cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register, cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in};

  //cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register <= 0;
      else 
        cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register <= p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
    end


  //local readdatavalid cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1, which is an e_mux
  assign cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1 = cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;

  assign cpu_2_data_master_requests_onchip_memory2_0_s1 = ({cpu_2_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h3000) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_onchip_memory2_0_s1 = cpu_2_data_master_requests_onchip_memory2_0_s1 & ~((cpu_2_data_master_read & ((1 < cpu_2_data_master_latency_counter) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in = cpu_2_data_master_granted_onchip_memory2_0_s1 & cpu_2_data_master_read & ~onchip_memory2_0_s1_waits_for_read;

  //shift register p1 cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register = {cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register, cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in};

  //cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register <= 0;
      else 
        cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register <= p1_cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
    end


  //local readdatavalid cpu_2_data_master_read_data_valid_onchip_memory2_0_s1, which is an e_mux
  assign cpu_2_data_master_read_data_valid_onchip_memory2_0_s1 = cpu_2_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;

  assign cpu_2_instruction_master_requests_onchip_memory2_0_s1 = (({cpu_2_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h3000) & (cpu_2_instruction_master_read)) & cpu_2_instruction_master_read;
  assign cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1 = cpu_2_instruction_master_requests_onchip_memory2_0_s1 & ~((cpu_2_instruction_master_read & ((1 < cpu_2_instruction_master_latency_counter) | (|cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in = cpu_2_instruction_master_granted_onchip_memory2_0_s1 & cpu_2_instruction_master_read & ~onchip_memory2_0_s1_waits_for_read;

  //shift register p1 cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register = {cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register, cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in};

  //cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register <= 0;
      else 
        cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register <= p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
    end


  //local readdatavalid cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1, which is an e_mux
  assign cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1 = cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;

  assign cpu_3_data_master_requests_onchip_memory2_0_s1 = ({cpu_3_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h3000) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_onchip_memory2_0_s1 = cpu_3_data_master_requests_onchip_memory2_0_s1 & ~((cpu_3_data_master_read & ((1 < cpu_3_data_master_latency_counter) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in = cpu_3_data_master_granted_onchip_memory2_0_s1 & cpu_3_data_master_read & ~onchip_memory2_0_s1_waits_for_read;

  //shift register p1 cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register = {cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register, cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register_in};

  //cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register <= 0;
      else 
        cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register <= p1_cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;
    end


  //local readdatavalid cpu_3_data_master_read_data_valid_onchip_memory2_0_s1, which is an e_mux
  assign cpu_3_data_master_read_data_valid_onchip_memory2_0_s1 = cpu_3_data_master_read_data_valid_onchip_memory2_0_s1_shift_register;

  assign cpu_3_instruction_master_requests_onchip_memory2_0_s1 = (({cpu_3_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h3000) & (cpu_3_instruction_master_read)) & cpu_3_instruction_master_read;
  assign cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1 = cpu_3_instruction_master_requests_onchip_memory2_0_s1 & ~((cpu_3_instruction_master_read & ((1 < cpu_3_instruction_master_latency_counter) | (|cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in = cpu_3_instruction_master_granted_onchip_memory2_0_s1 & cpu_3_instruction_master_read & ~onchip_memory2_0_s1_waits_for_read;

  //shift register p1 cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register = {cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register, cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register_in};

  //cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register <= 0;
      else 
        cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register <= p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;
    end


  //local readdatavalid cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1, which is an e_mux
  assign cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1 = cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1_shift_register;

  //allow new arb cycle for onchip_memory2_0/s1, which is an e_assign
  assign onchip_memory2_0_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_1_instruction_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_2_instruction_master_arbiterlock & ~cpu_3_data_master_arbiterlock & ~cpu_3_instruction_master_arbiterlock;

  //cpu_3/instruction_master assignment into master qualified-requests vector for onchip_memory2_0/s1, which is an e_assign
  assign onchip_memory2_0_s1_master_qreq_vector[0] = cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1;

  //cpu_3/instruction_master grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_3_instruction_master_granted_onchip_memory2_0_s1 = onchip_memory2_0_s1_grant_vector[0];

  //cpu_3/instruction_master saved-grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_3_instruction_master_saved_grant_onchip_memory2_0_s1 = onchip_memory2_0_s1_arb_winner[0] && cpu_3_instruction_master_requests_onchip_memory2_0_s1;

  //cpu_3/data_master assignment into master qualified-requests vector for onchip_memory2_0/s1, which is an e_assign
  assign onchip_memory2_0_s1_master_qreq_vector[1] = cpu_3_data_master_qualified_request_onchip_memory2_0_s1;

  //cpu_3/data_master grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_3_data_master_granted_onchip_memory2_0_s1 = onchip_memory2_0_s1_grant_vector[1];

  //cpu_3/data_master saved-grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_3_data_master_saved_grant_onchip_memory2_0_s1 = onchip_memory2_0_s1_arb_winner[1] && cpu_3_data_master_requests_onchip_memory2_0_s1;

  //cpu_2/instruction_master assignment into master qualified-requests vector for onchip_memory2_0/s1, which is an e_assign
  assign onchip_memory2_0_s1_master_qreq_vector[2] = cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1;

  //cpu_2/instruction_master grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_2_instruction_master_granted_onchip_memory2_0_s1 = onchip_memory2_0_s1_grant_vector[2];

  //cpu_2/instruction_master saved-grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_2_instruction_master_saved_grant_onchip_memory2_0_s1 = onchip_memory2_0_s1_arb_winner[2] && cpu_2_instruction_master_requests_onchip_memory2_0_s1;

  //cpu_2/data_master assignment into master qualified-requests vector for onchip_memory2_0/s1, which is an e_assign
  assign onchip_memory2_0_s1_master_qreq_vector[3] = cpu_2_data_master_qualified_request_onchip_memory2_0_s1;

  //cpu_2/data_master grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_2_data_master_granted_onchip_memory2_0_s1 = onchip_memory2_0_s1_grant_vector[3];

  //cpu_2/data_master saved-grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_2_data_master_saved_grant_onchip_memory2_0_s1 = onchip_memory2_0_s1_arb_winner[3] && cpu_2_data_master_requests_onchip_memory2_0_s1;

  //cpu_1/instruction_master assignment into master qualified-requests vector for onchip_memory2_0/s1, which is an e_assign
  assign onchip_memory2_0_s1_master_qreq_vector[4] = cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1;

  //cpu_1/instruction_master grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_1_instruction_master_granted_onchip_memory2_0_s1 = onchip_memory2_0_s1_grant_vector[4];

  //cpu_1/instruction_master saved-grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_1_instruction_master_saved_grant_onchip_memory2_0_s1 = onchip_memory2_0_s1_arb_winner[4] && cpu_1_instruction_master_requests_onchip_memory2_0_s1;

  //cpu_1/data_master assignment into master qualified-requests vector for onchip_memory2_0/s1, which is an e_assign
  assign onchip_memory2_0_s1_master_qreq_vector[5] = cpu_1_data_master_qualified_request_onchip_memory2_0_s1;

  //cpu_1/data_master grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_1_data_master_granted_onchip_memory2_0_s1 = onchip_memory2_0_s1_grant_vector[5];

  //cpu_1/data_master saved-grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_1_data_master_saved_grant_onchip_memory2_0_s1 = onchip_memory2_0_s1_arb_winner[5] && cpu_1_data_master_requests_onchip_memory2_0_s1;

  //cpu_0/instruction_master assignment into master qualified-requests vector for onchip_memory2_0/s1, which is an e_assign
  assign onchip_memory2_0_s1_master_qreq_vector[6] = cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1;

  //cpu_0/instruction_master grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_0_instruction_master_granted_onchip_memory2_0_s1 = onchip_memory2_0_s1_grant_vector[6];

  //cpu_0/instruction_master saved-grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_onchip_memory2_0_s1 = onchip_memory2_0_s1_arb_winner[6] && cpu_0_instruction_master_requests_onchip_memory2_0_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for onchip_memory2_0/s1, which is an e_assign
  assign onchip_memory2_0_s1_master_qreq_vector[7] = cpu_0_data_master_qualified_request_onchip_memory2_0_s1;

  //cpu_0/data_master grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_0_data_master_granted_onchip_memory2_0_s1 = onchip_memory2_0_s1_grant_vector[7];

  //cpu_0/data_master saved-grant onchip_memory2_0/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_onchip_memory2_0_s1 = onchip_memory2_0_s1_arb_winner[7] && cpu_0_data_master_requests_onchip_memory2_0_s1;

  //onchip_memory2_0/s1 chosen-master double-vector, which is an e_assign
  assign onchip_memory2_0_s1_chosen_master_double_vector = {onchip_memory2_0_s1_master_qreq_vector, onchip_memory2_0_s1_master_qreq_vector} & ({~onchip_memory2_0_s1_master_qreq_vector, ~onchip_memory2_0_s1_master_qreq_vector} + onchip_memory2_0_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign onchip_memory2_0_s1_arb_winner = (onchip_memory2_0_s1_allow_new_arb_cycle & | onchip_memory2_0_s1_grant_vector) ? onchip_memory2_0_s1_grant_vector : onchip_memory2_0_s1_saved_chosen_master_vector;

  //saved onchip_memory2_0_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_0_s1_saved_chosen_master_vector <= 0;
      else if (onchip_memory2_0_s1_allow_new_arb_cycle)
          onchip_memory2_0_s1_saved_chosen_master_vector <= |onchip_memory2_0_s1_grant_vector ? onchip_memory2_0_s1_grant_vector : onchip_memory2_0_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign onchip_memory2_0_s1_grant_vector = {(onchip_memory2_0_s1_chosen_master_double_vector[7] | onchip_memory2_0_s1_chosen_master_double_vector[15]),
    (onchip_memory2_0_s1_chosen_master_double_vector[6] | onchip_memory2_0_s1_chosen_master_double_vector[14]),
    (onchip_memory2_0_s1_chosen_master_double_vector[5] | onchip_memory2_0_s1_chosen_master_double_vector[13]),
    (onchip_memory2_0_s1_chosen_master_double_vector[4] | onchip_memory2_0_s1_chosen_master_double_vector[12]),
    (onchip_memory2_0_s1_chosen_master_double_vector[3] | onchip_memory2_0_s1_chosen_master_double_vector[11]),
    (onchip_memory2_0_s1_chosen_master_double_vector[2] | onchip_memory2_0_s1_chosen_master_double_vector[10]),
    (onchip_memory2_0_s1_chosen_master_double_vector[1] | onchip_memory2_0_s1_chosen_master_double_vector[9]),
    (onchip_memory2_0_s1_chosen_master_double_vector[0] | onchip_memory2_0_s1_chosen_master_double_vector[8])};

  //onchip_memory2_0/s1 chosen master rotated left, which is an e_assign
  assign onchip_memory2_0_s1_chosen_master_rot_left = (onchip_memory2_0_s1_arb_winner << 1) ? (onchip_memory2_0_s1_arb_winner << 1) : 1;

  //onchip_memory2_0/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_0_s1_arb_addend <= 1;
      else if (|onchip_memory2_0_s1_grant_vector)
          onchip_memory2_0_s1_arb_addend <= onchip_memory2_0_s1_end_xfer? onchip_memory2_0_s1_chosen_master_rot_left : onchip_memory2_0_s1_grant_vector;
    end


  //~onchip_memory2_0_s1_reset assignment, which is an e_assign
  assign onchip_memory2_0_s1_reset = ~reset_n;

  assign onchip_memory2_0_s1_chipselect = cpu_0_data_master_granted_onchip_memory2_0_s1 | cpu_0_instruction_master_granted_onchip_memory2_0_s1 | cpu_1_data_master_granted_onchip_memory2_0_s1 | cpu_1_instruction_master_granted_onchip_memory2_0_s1 | cpu_2_data_master_granted_onchip_memory2_0_s1 | cpu_2_instruction_master_granted_onchip_memory2_0_s1 | cpu_3_data_master_granted_onchip_memory2_0_s1 | cpu_3_instruction_master_granted_onchip_memory2_0_s1;
  //onchip_memory2_0_s1_firsttransfer first transaction, which is an e_assign
  assign onchip_memory2_0_s1_firsttransfer = onchip_memory2_0_s1_begins_xfer ? onchip_memory2_0_s1_unreg_firsttransfer : onchip_memory2_0_s1_reg_firsttransfer;

  //onchip_memory2_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign onchip_memory2_0_s1_unreg_firsttransfer = ~(onchip_memory2_0_s1_slavearbiterlockenable & onchip_memory2_0_s1_any_continuerequest);

  //onchip_memory2_0_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_0_s1_reg_firsttransfer <= 1'b1;
      else if (onchip_memory2_0_s1_begins_xfer)
          onchip_memory2_0_s1_reg_firsttransfer <= onchip_memory2_0_s1_unreg_firsttransfer;
    end


  //onchip_memory2_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign onchip_memory2_0_s1_beginbursttransfer_internal = onchip_memory2_0_s1_begins_xfer;

  //onchip_memory2_0_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign onchip_memory2_0_s1_arbitration_holdoff_internal = onchip_memory2_0_s1_begins_xfer & onchip_memory2_0_s1_firsttransfer;

  //onchip_memory2_0_s1_write assignment, which is an e_mux
  assign onchip_memory2_0_s1_write = (cpu_0_data_master_granted_onchip_memory2_0_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_onchip_memory2_0_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_onchip_memory2_0_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_onchip_memory2_0_s1 & cpu_3_data_master_write);

  assign shifted_address_to_onchip_memory2_0_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //onchip_memory2_0_s1_address mux, which is an e_mux
  assign onchip_memory2_0_s1_address = (cpu_0_data_master_granted_onchip_memory2_0_s1)? (shifted_address_to_onchip_memory2_0_s1_from_cpu_0_data_master >> 2) :
    (cpu_0_instruction_master_granted_onchip_memory2_0_s1)? (shifted_address_to_onchip_memory2_0_s1_from_cpu_0_instruction_master >> 2) :
    (cpu_1_data_master_granted_onchip_memory2_0_s1)? (shifted_address_to_onchip_memory2_0_s1_from_cpu_1_data_master >> 2) :
    (cpu_1_instruction_master_granted_onchip_memory2_0_s1)? (shifted_address_to_onchip_memory2_0_s1_from_cpu_1_instruction_master >> 2) :
    (cpu_2_data_master_granted_onchip_memory2_0_s1)? (shifted_address_to_onchip_memory2_0_s1_from_cpu_2_data_master >> 2) :
    (cpu_2_instruction_master_granted_onchip_memory2_0_s1)? (shifted_address_to_onchip_memory2_0_s1_from_cpu_2_instruction_master >> 2) :
    (cpu_3_data_master_granted_onchip_memory2_0_s1)? (shifted_address_to_onchip_memory2_0_s1_from_cpu_3_data_master >> 2) :
    (shifted_address_to_onchip_memory2_0_s1_from_cpu_3_instruction_master >> 2);

  assign shifted_address_to_onchip_memory2_0_s1_from_cpu_0_instruction_master = cpu_0_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_0_s1_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_0_s1_from_cpu_1_instruction_master = cpu_1_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_0_s1_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_0_s1_from_cpu_2_instruction_master = cpu_2_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_0_s1_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_0_s1_from_cpu_3_instruction_master = cpu_3_instruction_master_address_to_slave;
  //d1_onchip_memory2_0_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_onchip_memory2_0_s1_end_xfer <= 1;
      else 
        d1_onchip_memory2_0_s1_end_xfer <= onchip_memory2_0_s1_end_xfer;
    end


  //onchip_memory2_0_s1_waits_for_read in a cycle, which is an e_mux
  assign onchip_memory2_0_s1_waits_for_read = onchip_memory2_0_s1_in_a_read_cycle & 0;

  //onchip_memory2_0_s1_in_a_read_cycle assignment, which is an e_assign
  assign onchip_memory2_0_s1_in_a_read_cycle = (cpu_0_data_master_granted_onchip_memory2_0_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_onchip_memory2_0_s1 & cpu_0_instruction_master_read) | (cpu_1_data_master_granted_onchip_memory2_0_s1 & cpu_1_data_master_read) | (cpu_1_instruction_master_granted_onchip_memory2_0_s1 & cpu_1_instruction_master_read) | (cpu_2_data_master_granted_onchip_memory2_0_s1 & cpu_2_data_master_read) | (cpu_2_instruction_master_granted_onchip_memory2_0_s1 & cpu_2_instruction_master_read) | (cpu_3_data_master_granted_onchip_memory2_0_s1 & cpu_3_data_master_read) | (cpu_3_instruction_master_granted_onchip_memory2_0_s1 & cpu_3_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = onchip_memory2_0_s1_in_a_read_cycle;

  //onchip_memory2_0_s1_waits_for_write in a cycle, which is an e_mux
  assign onchip_memory2_0_s1_waits_for_write = onchip_memory2_0_s1_in_a_write_cycle & 0;

  //onchip_memory2_0_s1_in_a_write_cycle assignment, which is an e_assign
  assign onchip_memory2_0_s1_in_a_write_cycle = (cpu_0_data_master_granted_onchip_memory2_0_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_onchip_memory2_0_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_onchip_memory2_0_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_onchip_memory2_0_s1 & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = onchip_memory2_0_s1_in_a_write_cycle;

  assign wait_for_onchip_memory2_0_s1_counter = 0;
  //onchip_memory2_0_s1_byteenable byte enable port mux, which is an e_mux
  assign onchip_memory2_0_s1_byteenable = (cpu_0_data_master_granted_onchip_memory2_0_s1)? cpu_0_data_master_byteenable :
    (cpu_1_data_master_granted_onchip_memory2_0_s1)? cpu_1_data_master_byteenable :
    (cpu_2_data_master_granted_onchip_memory2_0_s1)? cpu_2_data_master_byteenable :
    (cpu_3_data_master_granted_onchip_memory2_0_s1)? cpu_3_data_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //onchip_memory2_0/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_onchip_memory2_0_s1 + cpu_0_instruction_master_granted_onchip_memory2_0_s1 + cpu_1_data_master_granted_onchip_memory2_0_s1 + cpu_1_instruction_master_granted_onchip_memory2_0_s1 + cpu_2_data_master_granted_onchip_memory2_0_s1 + cpu_2_instruction_master_granted_onchip_memory2_0_s1 + cpu_3_data_master_granted_onchip_memory2_0_s1 + cpu_3_instruction_master_granted_onchip_memory2_0_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_onchip_memory2_0_s1 + cpu_0_instruction_master_saved_grant_onchip_memory2_0_s1 + cpu_1_data_master_saved_grant_onchip_memory2_0_s1 + cpu_1_instruction_master_saved_grant_onchip_memory2_0_s1 + cpu_2_data_master_saved_grant_onchip_memory2_0_s1 + cpu_2_instruction_master_saved_grant_onchip_memory2_0_s1 + cpu_3_data_master_saved_grant_onchip_memory2_0_s1 + cpu_3_instruction_master_saved_grant_onchip_memory2_0_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module onchip_memory2_1_s1_arbitrator (
                                        // inputs:
                                         clk,
                                         cpu_0_data_master_address_to_slave,
                                         cpu_0_data_master_byteenable,
                                         cpu_0_data_master_latency_counter,
                                         cpu_0_data_master_read,
                                         cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_0_data_master_write,
                                         cpu_0_data_master_writedata,
                                         cpu_0_instruction_master_address_to_slave,
                                         cpu_0_instruction_master_latency_counter,
                                         cpu_0_instruction_master_read,
                                         cpu_1_data_master_address_to_slave,
                                         cpu_1_data_master_byteenable,
                                         cpu_1_data_master_latency_counter,
                                         cpu_1_data_master_read,
                                         cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_1_data_master_write,
                                         cpu_1_data_master_writedata,
                                         cpu_1_instruction_master_address_to_slave,
                                         cpu_1_instruction_master_latency_counter,
                                         cpu_1_instruction_master_read,
                                         cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_2_data_master_address_to_slave,
                                         cpu_2_data_master_byteenable,
                                         cpu_2_data_master_latency_counter,
                                         cpu_2_data_master_read,
                                         cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_2_data_master_write,
                                         cpu_2_data_master_writedata,
                                         cpu_2_instruction_master_address_to_slave,
                                         cpu_2_instruction_master_latency_counter,
                                         cpu_2_instruction_master_read,
                                         cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_3_data_master_address_to_slave,
                                         cpu_3_data_master_byteenable,
                                         cpu_3_data_master_latency_counter,
                                         cpu_3_data_master_read,
                                         cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_3_data_master_write,
                                         cpu_3_data_master_writedata,
                                         cpu_3_instruction_master_address_to_slave,
                                         cpu_3_instruction_master_latency_counter,
                                         cpu_3_instruction_master_read,
                                         cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         onchip_memory2_1_s1_readdata,
                                         reset_n,

                                        // outputs:
                                         cpu_0_data_master_granted_onchip_memory2_1_s1,
                                         cpu_0_data_master_qualified_request_onchip_memory2_1_s1,
                                         cpu_0_data_master_read_data_valid_onchip_memory2_1_s1,
                                         cpu_0_data_master_requests_onchip_memory2_1_s1,
                                         cpu_0_instruction_master_granted_onchip_memory2_1_s1,
                                         cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1,
                                         cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1,
                                         cpu_0_instruction_master_requests_onchip_memory2_1_s1,
                                         cpu_1_data_master_granted_onchip_memory2_1_s1,
                                         cpu_1_data_master_qualified_request_onchip_memory2_1_s1,
                                         cpu_1_data_master_read_data_valid_onchip_memory2_1_s1,
                                         cpu_1_data_master_requests_onchip_memory2_1_s1,
                                         cpu_1_instruction_master_granted_onchip_memory2_1_s1,
                                         cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1,
                                         cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1,
                                         cpu_1_instruction_master_requests_onchip_memory2_1_s1,
                                         cpu_2_data_master_granted_onchip_memory2_1_s1,
                                         cpu_2_data_master_qualified_request_onchip_memory2_1_s1,
                                         cpu_2_data_master_read_data_valid_onchip_memory2_1_s1,
                                         cpu_2_data_master_requests_onchip_memory2_1_s1,
                                         cpu_2_instruction_master_granted_onchip_memory2_1_s1,
                                         cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1,
                                         cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1,
                                         cpu_2_instruction_master_requests_onchip_memory2_1_s1,
                                         cpu_3_data_master_granted_onchip_memory2_1_s1,
                                         cpu_3_data_master_qualified_request_onchip_memory2_1_s1,
                                         cpu_3_data_master_read_data_valid_onchip_memory2_1_s1,
                                         cpu_3_data_master_requests_onchip_memory2_1_s1,
                                         cpu_3_instruction_master_granted_onchip_memory2_1_s1,
                                         cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1,
                                         cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1,
                                         cpu_3_instruction_master_requests_onchip_memory2_1_s1,
                                         d1_onchip_memory2_1_s1_end_xfer,
                                         onchip_memory2_1_s1_address,
                                         onchip_memory2_1_s1_byteenable,
                                         onchip_memory2_1_s1_chipselect,
                                         onchip_memory2_1_s1_clken,
                                         onchip_memory2_1_s1_readdata_from_sa,
                                         onchip_memory2_1_s1_reset,
                                         onchip_memory2_1_s1_write,
                                         onchip_memory2_1_s1_writedata
                                      )
;

  output           cpu_0_data_master_granted_onchip_memory2_1_s1;
  output           cpu_0_data_master_qualified_request_onchip_memory2_1_s1;
  output           cpu_0_data_master_read_data_valid_onchip_memory2_1_s1;
  output           cpu_0_data_master_requests_onchip_memory2_1_s1;
  output           cpu_0_instruction_master_granted_onchip_memory2_1_s1;
  output           cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1;
  output           cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1;
  output           cpu_0_instruction_master_requests_onchip_memory2_1_s1;
  output           cpu_1_data_master_granted_onchip_memory2_1_s1;
  output           cpu_1_data_master_qualified_request_onchip_memory2_1_s1;
  output           cpu_1_data_master_read_data_valid_onchip_memory2_1_s1;
  output           cpu_1_data_master_requests_onchip_memory2_1_s1;
  output           cpu_1_instruction_master_granted_onchip_memory2_1_s1;
  output           cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1;
  output           cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1;
  output           cpu_1_instruction_master_requests_onchip_memory2_1_s1;
  output           cpu_2_data_master_granted_onchip_memory2_1_s1;
  output           cpu_2_data_master_qualified_request_onchip_memory2_1_s1;
  output           cpu_2_data_master_read_data_valid_onchip_memory2_1_s1;
  output           cpu_2_data_master_requests_onchip_memory2_1_s1;
  output           cpu_2_instruction_master_granted_onchip_memory2_1_s1;
  output           cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1;
  output           cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1;
  output           cpu_2_instruction_master_requests_onchip_memory2_1_s1;
  output           cpu_3_data_master_granted_onchip_memory2_1_s1;
  output           cpu_3_data_master_qualified_request_onchip_memory2_1_s1;
  output           cpu_3_data_master_read_data_valid_onchip_memory2_1_s1;
  output           cpu_3_data_master_requests_onchip_memory2_1_s1;
  output           cpu_3_instruction_master_granted_onchip_memory2_1_s1;
  output           cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1;
  output           cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1;
  output           cpu_3_instruction_master_requests_onchip_memory2_1_s1;
  output           d1_onchip_memory2_1_s1_end_xfer;
  output  [  6: 0] onchip_memory2_1_s1_address;
  output  [  3: 0] onchip_memory2_1_s1_byteenable;
  output           onchip_memory2_1_s1_chipselect;
  output           onchip_memory2_1_s1_clken;
  output  [ 31: 0] onchip_memory2_1_s1_readdata_from_sa;
  output           onchip_memory2_1_s1_reset;
  output           onchip_memory2_1_s1_write;
  output  [ 31: 0] onchip_memory2_1_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input            cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input   [  3: 0] cpu_1_data_master_byteenable;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_1_instruction_master_address_to_slave;
  input            cpu_1_instruction_master_latency_counter;
  input            cpu_1_instruction_master_read;
  input            cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input   [  3: 0] cpu_2_data_master_byteenable;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_2_instruction_master_address_to_slave;
  input            cpu_2_instruction_master_latency_counter;
  input            cpu_2_instruction_master_read;
  input            cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input   [  3: 0] cpu_3_data_master_byteenable;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 24: 0] cpu_3_instruction_master_address_to_slave;
  input            cpu_3_instruction_master_latency_counter;
  input            cpu_3_instruction_master_read;
  input            cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 31: 0] onchip_memory2_1_s1_readdata;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_onchip_memory2_1_s1;
  wire             cpu_0_data_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_1_s1;
  reg              cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in;
  wire             cpu_0_data_master_requests_onchip_memory2_1_s1;
  wire             cpu_0_data_master_saved_grant_onchip_memory2_1_s1;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_onchip_memory2_1_s1;
  wire             cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1;
  reg              cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in;
  wire             cpu_0_instruction_master_requests_onchip_memory2_1_s1;
  wire             cpu_0_instruction_master_saved_grant_onchip_memory2_1_s1;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_onchip_memory2_1_s1;
  wire             cpu_1_data_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_1_s1;
  reg              cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in;
  wire             cpu_1_data_master_requests_onchip_memory2_1_s1;
  wire             cpu_1_data_master_saved_grant_onchip_memory2_1_s1;
  wire             cpu_1_instruction_master_arbiterlock;
  wire             cpu_1_instruction_master_arbiterlock2;
  wire             cpu_1_instruction_master_continuerequest;
  wire             cpu_1_instruction_master_granted_onchip_memory2_1_s1;
  wire             cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1;
  reg              cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in;
  wire             cpu_1_instruction_master_requests_onchip_memory2_1_s1;
  wire             cpu_1_instruction_master_saved_grant_onchip_memory2_1_s1;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_onchip_memory2_1_s1;
  wire             cpu_2_data_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_1_s1;
  reg              cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in;
  wire             cpu_2_data_master_requests_onchip_memory2_1_s1;
  wire             cpu_2_data_master_saved_grant_onchip_memory2_1_s1;
  wire             cpu_2_instruction_master_arbiterlock;
  wire             cpu_2_instruction_master_arbiterlock2;
  wire             cpu_2_instruction_master_continuerequest;
  wire             cpu_2_instruction_master_granted_onchip_memory2_1_s1;
  wire             cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1;
  reg              cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in;
  wire             cpu_2_instruction_master_requests_onchip_memory2_1_s1;
  wire             cpu_2_instruction_master_saved_grant_onchip_memory2_1_s1;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_onchip_memory2_1_s1;
  wire             cpu_3_data_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_1_s1;
  reg              cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in;
  wire             cpu_3_data_master_requests_onchip_memory2_1_s1;
  wire             cpu_3_data_master_saved_grant_onchip_memory2_1_s1;
  wire             cpu_3_instruction_master_arbiterlock;
  wire             cpu_3_instruction_master_arbiterlock2;
  wire             cpu_3_instruction_master_continuerequest;
  wire             cpu_3_instruction_master_granted_onchip_memory2_1_s1;
  wire             cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1;
  reg              cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in;
  wire             cpu_3_instruction_master_requests_onchip_memory2_1_s1;
  wire             cpu_3_instruction_master_saved_grant_onchip_memory2_1_s1;
  reg              d1_onchip_memory2_1_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_onchip_memory2_1_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_1_s1;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_1_s1;
  reg              last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_1_s1;
  reg              last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_1_s1;
  reg              last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_1_s1;
  reg              last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_1_s1;
  reg              last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_1_s1;
  reg              last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_1_s1;
  wire    [  6: 0] onchip_memory2_1_s1_address;
  wire             onchip_memory2_1_s1_allgrants;
  wire             onchip_memory2_1_s1_allow_new_arb_cycle;
  wire             onchip_memory2_1_s1_any_bursting_master_saved_grant;
  wire             onchip_memory2_1_s1_any_continuerequest;
  reg     [  7: 0] onchip_memory2_1_s1_arb_addend;
  wire             onchip_memory2_1_s1_arb_counter_enable;
  reg     [  2: 0] onchip_memory2_1_s1_arb_share_counter;
  wire    [  2: 0] onchip_memory2_1_s1_arb_share_counter_next_value;
  wire    [  2: 0] onchip_memory2_1_s1_arb_share_set_values;
  wire    [  7: 0] onchip_memory2_1_s1_arb_winner;
  wire             onchip_memory2_1_s1_arbitration_holdoff_internal;
  wire             onchip_memory2_1_s1_beginbursttransfer_internal;
  wire             onchip_memory2_1_s1_begins_xfer;
  wire    [  3: 0] onchip_memory2_1_s1_byteenable;
  wire             onchip_memory2_1_s1_chipselect;
  wire    [ 15: 0] onchip_memory2_1_s1_chosen_master_double_vector;
  wire    [  7: 0] onchip_memory2_1_s1_chosen_master_rot_left;
  wire             onchip_memory2_1_s1_clken;
  wire             onchip_memory2_1_s1_end_xfer;
  wire             onchip_memory2_1_s1_firsttransfer;
  wire    [  7: 0] onchip_memory2_1_s1_grant_vector;
  wire             onchip_memory2_1_s1_in_a_read_cycle;
  wire             onchip_memory2_1_s1_in_a_write_cycle;
  wire    [  7: 0] onchip_memory2_1_s1_master_qreq_vector;
  wire             onchip_memory2_1_s1_non_bursting_master_requests;
  wire    [ 31: 0] onchip_memory2_1_s1_readdata_from_sa;
  reg              onchip_memory2_1_s1_reg_firsttransfer;
  wire             onchip_memory2_1_s1_reset;
  reg     [  7: 0] onchip_memory2_1_s1_saved_chosen_master_vector;
  reg              onchip_memory2_1_s1_slavearbiterlockenable;
  wire             onchip_memory2_1_s1_slavearbiterlockenable2;
  wire             onchip_memory2_1_s1_unreg_firsttransfer;
  wire             onchip_memory2_1_s1_waits_for_read;
  wire             onchip_memory2_1_s1_waits_for_write;
  wire             onchip_memory2_1_s1_write;
  wire    [ 31: 0] onchip_memory2_1_s1_writedata;
  wire             p1_cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             p1_cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             p1_cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             p1_cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire             p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_1_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_1_s1_from_cpu_0_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_1_s1_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_1_s1_from_cpu_1_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_1_s1_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_1_s1_from_cpu_2_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_1_s1_from_cpu_3_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_1_s1_from_cpu_3_instruction_master;
  wire             wait_for_onchip_memory2_1_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~onchip_memory2_1_s1_end_xfer;
    end


  assign onchip_memory2_1_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_onchip_memory2_1_s1 | cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1 | cpu_1_data_master_qualified_request_onchip_memory2_1_s1 | cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1 | cpu_2_data_master_qualified_request_onchip_memory2_1_s1 | cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1 | cpu_3_data_master_qualified_request_onchip_memory2_1_s1 | cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1));
  //assign onchip_memory2_1_s1_readdata_from_sa = onchip_memory2_1_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign onchip_memory2_1_s1_readdata_from_sa = onchip_memory2_1_s1_readdata;

  assign cpu_0_data_master_requests_onchip_memory2_1_s1 = ({cpu_0_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h4000) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //onchip_memory2_1_s1_arb_share_counter set values, which is an e_mux
  assign onchip_memory2_1_s1_arb_share_set_values = 1;

  //onchip_memory2_1_s1_non_bursting_master_requests mux, which is an e_mux
  assign onchip_memory2_1_s1_non_bursting_master_requests = cpu_0_data_master_requests_onchip_memory2_1_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_1_data_master_requests_onchip_memory2_1_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_2_data_master_requests_onchip_memory2_1_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_3_data_master_requests_onchip_memory2_1_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_0_data_master_requests_onchip_memory2_1_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_1_data_master_requests_onchip_memory2_1_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_2_data_master_requests_onchip_memory2_1_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_3_data_master_requests_onchip_memory2_1_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_0_data_master_requests_onchip_memory2_1_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_1_data_master_requests_onchip_memory2_1_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_2_data_master_requests_onchip_memory2_1_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_3_data_master_requests_onchip_memory2_1_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_0_data_master_requests_onchip_memory2_1_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_1_data_master_requests_onchip_memory2_1_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_2_data_master_requests_onchip_memory2_1_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_3_data_master_requests_onchip_memory2_1_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_0_data_master_requests_onchip_memory2_1_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_1_data_master_requests_onchip_memory2_1_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_2_data_master_requests_onchip_memory2_1_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_3_data_master_requests_onchip_memory2_1_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_0_data_master_requests_onchip_memory2_1_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_1_data_master_requests_onchip_memory2_1_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_2_data_master_requests_onchip_memory2_1_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_3_data_master_requests_onchip_memory2_1_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_0_data_master_requests_onchip_memory2_1_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_1_data_master_requests_onchip_memory2_1_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_2_data_master_requests_onchip_memory2_1_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_3_data_master_requests_onchip_memory2_1_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_0_data_master_requests_onchip_memory2_1_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_1_data_master_requests_onchip_memory2_1_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_2_data_master_requests_onchip_memory2_1_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_1_s1 |
    cpu_3_data_master_requests_onchip_memory2_1_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_1_s1;

  //onchip_memory2_1_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign onchip_memory2_1_s1_any_bursting_master_saved_grant = 0;

  //onchip_memory2_1_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign onchip_memory2_1_s1_arb_share_counter_next_value = onchip_memory2_1_s1_firsttransfer ? (onchip_memory2_1_s1_arb_share_set_values - 1) : |onchip_memory2_1_s1_arb_share_counter ? (onchip_memory2_1_s1_arb_share_counter - 1) : 0;

  //onchip_memory2_1_s1_allgrants all slave grants, which is an e_mux
  assign onchip_memory2_1_s1_allgrants = (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector) |
    (|onchip_memory2_1_s1_grant_vector);

  //onchip_memory2_1_s1_end_xfer assignment, which is an e_assign
  assign onchip_memory2_1_s1_end_xfer = ~(onchip_memory2_1_s1_waits_for_read | onchip_memory2_1_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_onchip_memory2_1_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_onchip_memory2_1_s1 = onchip_memory2_1_s1_end_xfer & (~onchip_memory2_1_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //onchip_memory2_1_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign onchip_memory2_1_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_onchip_memory2_1_s1 & onchip_memory2_1_s1_allgrants) | (end_xfer_arb_share_counter_term_onchip_memory2_1_s1 & ~onchip_memory2_1_s1_non_bursting_master_requests);

  //onchip_memory2_1_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_1_s1_arb_share_counter <= 0;
      else if (onchip_memory2_1_s1_arb_counter_enable)
          onchip_memory2_1_s1_arb_share_counter <= onchip_memory2_1_s1_arb_share_counter_next_value;
    end


  //onchip_memory2_1_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_1_s1_slavearbiterlockenable <= 0;
      else if ((|onchip_memory2_1_s1_master_qreq_vector & end_xfer_arb_share_counter_term_onchip_memory2_1_s1) | (end_xfer_arb_share_counter_term_onchip_memory2_1_s1 & ~onchip_memory2_1_s1_non_bursting_master_requests))
          onchip_memory2_1_s1_slavearbiterlockenable <= |onchip_memory2_1_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master onchip_memory2_1/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = onchip_memory2_1_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //onchip_memory2_1_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign onchip_memory2_1_s1_slavearbiterlockenable2 = |onchip_memory2_1_s1_arb_share_counter_next_value;

  //cpu_0/data_master onchip_memory2_1/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = onchip_memory2_1_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master onchip_memory2_1/s1 arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = onchip_memory2_1_s1_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master onchip_memory2_1/s1 arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = onchip_memory2_1_s1_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted onchip_memory2_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_1_s1 <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_1_s1 <= cpu_0_instruction_master_saved_grant_onchip_memory2_1_s1 ? 1 : (onchip_memory2_1_s1_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_onchip_memory2_1_s1) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_1_s1;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_0_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_0_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_0_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_0_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_0_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_0_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_0_instruction_master_requests_onchip_memory2_1_s1);

  //onchip_memory2_1_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign onchip_memory2_1_s1_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest;

  //cpu_1/data_master onchip_memory2_1/s1 arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = onchip_memory2_1_s1_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master onchip_memory2_1/s1 arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = onchip_memory2_1_s1_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted onchip_memory2_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_1_s1 <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_1_s1 <= cpu_1_data_master_saved_grant_onchip_memory2_1_s1 ? 1 : (onchip_memory2_1_s1_arbitration_holdoff_internal | ~cpu_1_data_master_requests_onchip_memory2_1_s1) ? 0 : last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_1_s1;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_1_s1 & cpu_1_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_1_s1 & cpu_1_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_1_s1 & cpu_1_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_1_s1 & cpu_1_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_1_s1 & cpu_1_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_1_s1 & cpu_1_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_1_s1 & cpu_1_data_master_requests_onchip_memory2_1_s1);

  //cpu_1/instruction_master onchip_memory2_1/s1 arbiterlock, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock = onchip_memory2_1_s1_slavearbiterlockenable & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master onchip_memory2_1/s1 arbiterlock2, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock2 = onchip_memory2_1_s1_slavearbiterlockenable2 & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master granted onchip_memory2_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_1_s1 <= 0;
      else 
        last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_1_s1 <= cpu_1_instruction_master_saved_grant_onchip_memory2_1_s1 ? 1 : (onchip_memory2_1_s1_arbitration_holdoff_internal | ~cpu_1_instruction_master_requests_onchip_memory2_1_s1) ? 0 : last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_1_s1;
    end


  //cpu_1_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_1_instruction_master_continuerequest = (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_1_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_1_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_1_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_1_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_1_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_1_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_1_instruction_master_requests_onchip_memory2_1_s1);

  //cpu_2/data_master onchip_memory2_1/s1 arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = onchip_memory2_1_s1_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master onchip_memory2_1/s1 arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = onchip_memory2_1_s1_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted onchip_memory2_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_1_s1 <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_1_s1 <= cpu_2_data_master_saved_grant_onchip_memory2_1_s1 ? 1 : (onchip_memory2_1_s1_arbitration_holdoff_internal | ~cpu_2_data_master_requests_onchip_memory2_1_s1) ? 0 : last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_1_s1;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_1_s1 & cpu_2_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_1_s1 & cpu_2_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_1_s1 & cpu_2_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_1_s1 & cpu_2_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_1_s1 & cpu_2_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_1_s1 & cpu_2_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_1_s1 & cpu_2_data_master_requests_onchip_memory2_1_s1);

  //cpu_2/instruction_master onchip_memory2_1/s1 arbiterlock, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock = onchip_memory2_1_s1_slavearbiterlockenable & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master onchip_memory2_1/s1 arbiterlock2, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock2 = onchip_memory2_1_s1_slavearbiterlockenable2 & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master granted onchip_memory2_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_1_s1 <= 0;
      else 
        last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_1_s1 <= cpu_2_instruction_master_saved_grant_onchip_memory2_1_s1 ? 1 : (onchip_memory2_1_s1_arbitration_holdoff_internal | ~cpu_2_instruction_master_requests_onchip_memory2_1_s1) ? 0 : last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_1_s1;
    end


  //cpu_2_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_2_instruction_master_continuerequest = (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_2_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_2_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_2_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_2_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_2_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_2_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_2_instruction_master_requests_onchip_memory2_1_s1);

  //cpu_3/data_master onchip_memory2_1/s1 arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = onchip_memory2_1_s1_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master onchip_memory2_1/s1 arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = onchip_memory2_1_s1_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted onchip_memory2_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_1_s1 <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_1_s1 <= cpu_3_data_master_saved_grant_onchip_memory2_1_s1 ? 1 : (onchip_memory2_1_s1_arbitration_holdoff_internal | ~cpu_3_data_master_requests_onchip_memory2_1_s1) ? 0 : last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_1_s1;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_1_s1 & cpu_3_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_1_s1 & cpu_3_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_1_s1 & cpu_3_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_1_s1 & cpu_3_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_1_s1 & cpu_3_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_1_s1 & cpu_3_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_1_s1 & cpu_3_data_master_requests_onchip_memory2_1_s1);

  //cpu_3/instruction_master onchip_memory2_1/s1 arbiterlock, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock = onchip_memory2_1_s1_slavearbiterlockenable & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master onchip_memory2_1/s1 arbiterlock2, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock2 = onchip_memory2_1_s1_slavearbiterlockenable2 & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master granted onchip_memory2_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_1_s1 <= 0;
      else 
        last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_1_s1 <= cpu_3_instruction_master_saved_grant_onchip_memory2_1_s1 ? 1 : (onchip_memory2_1_s1_arbitration_holdoff_internal | ~cpu_3_instruction_master_requests_onchip_memory2_1_s1) ? 0 : last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_1_s1;
    end


  //cpu_3_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_3_instruction_master_continuerequest = (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_3_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_3_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_3_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_3_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_3_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_3_instruction_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_1_s1 & cpu_3_instruction_master_requests_onchip_memory2_1_s1);

  assign cpu_0_data_master_qualified_request_onchip_memory2_1_s1 = cpu_0_data_master_requests_onchip_memory2_1_s1 & ~((cpu_0_data_master_read & ((1 < cpu_0_data_master_latency_counter) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in = cpu_0_data_master_granted_onchip_memory2_1_s1 & cpu_0_data_master_read & ~onchip_memory2_1_s1_waits_for_read;

  //shift register p1 cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register = {cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register, cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in};

  //cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register <= 0;
      else 
        cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register <= p1_cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
    end


  //local readdatavalid cpu_0_data_master_read_data_valid_onchip_memory2_1_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_onchip_memory2_1_s1 = cpu_0_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;

  //onchip_memory2_1_s1_writedata mux, which is an e_mux
  assign onchip_memory2_1_s1_writedata = (cpu_0_data_master_granted_onchip_memory2_1_s1)? cpu_0_data_master_writedata :
    (cpu_1_data_master_granted_onchip_memory2_1_s1)? cpu_1_data_master_writedata :
    (cpu_2_data_master_granted_onchip_memory2_1_s1)? cpu_2_data_master_writedata :
    cpu_3_data_master_writedata;

  //mux onchip_memory2_1_s1_clken, which is an e_mux
  assign onchip_memory2_1_s1_clken = 1'b1;

  assign cpu_0_instruction_master_requests_onchip_memory2_1_s1 = (({cpu_0_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h4000) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted onchip_memory2_1/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_1_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_1_s1 <= cpu_0_data_master_saved_grant_onchip_memory2_1_s1 ? 1 : (onchip_memory2_1_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_onchip_memory2_1_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_1_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_1_s1 & cpu_0_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_1_s1 & cpu_0_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_1_s1 & cpu_0_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_1_s1 & cpu_0_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_1_s1 & cpu_0_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_1_s1 & cpu_0_data_master_requests_onchip_memory2_1_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_1_s1 & cpu_0_data_master_requests_onchip_memory2_1_s1);

  assign cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1 = cpu_0_instruction_master_requests_onchip_memory2_1_s1 & ~((cpu_0_instruction_master_read & ((1 < cpu_0_instruction_master_latency_counter))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in = cpu_0_instruction_master_granted_onchip_memory2_1_s1 & cpu_0_instruction_master_read & ~onchip_memory2_1_s1_waits_for_read;

  //shift register p1 cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register = {cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register, cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in};

  //cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register <= 0;
      else 
        cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register <= p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
    end


  //local readdatavalid cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1 = cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;

  assign cpu_1_data_master_requests_onchip_memory2_1_s1 = ({cpu_1_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h4000) & (cpu_1_data_master_read | cpu_1_data_master_write);
  assign cpu_1_data_master_qualified_request_onchip_memory2_1_s1 = cpu_1_data_master_requests_onchip_memory2_1_s1 & ~((cpu_1_data_master_read & ((1 < cpu_1_data_master_latency_counter) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in = cpu_1_data_master_granted_onchip_memory2_1_s1 & cpu_1_data_master_read & ~onchip_memory2_1_s1_waits_for_read;

  //shift register p1 cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register = {cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register, cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in};

  //cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register <= 0;
      else 
        cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register <= p1_cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
    end


  //local readdatavalid cpu_1_data_master_read_data_valid_onchip_memory2_1_s1, which is an e_mux
  assign cpu_1_data_master_read_data_valid_onchip_memory2_1_s1 = cpu_1_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;

  assign cpu_1_instruction_master_requests_onchip_memory2_1_s1 = (({cpu_1_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h4000) & (cpu_1_instruction_master_read)) & cpu_1_instruction_master_read;
  assign cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1 = cpu_1_instruction_master_requests_onchip_memory2_1_s1 & ~((cpu_1_instruction_master_read & ((1 < cpu_1_instruction_master_latency_counter) | (|cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in = cpu_1_instruction_master_granted_onchip_memory2_1_s1 & cpu_1_instruction_master_read & ~onchip_memory2_1_s1_waits_for_read;

  //shift register p1 cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register = {cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register, cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in};

  //cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register <= 0;
      else 
        cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register <= p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
    end


  //local readdatavalid cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1, which is an e_mux
  assign cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1 = cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;

  assign cpu_2_data_master_requests_onchip_memory2_1_s1 = ({cpu_2_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h4000) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_onchip_memory2_1_s1 = cpu_2_data_master_requests_onchip_memory2_1_s1 & ~((cpu_2_data_master_read & ((1 < cpu_2_data_master_latency_counter) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in = cpu_2_data_master_granted_onchip_memory2_1_s1 & cpu_2_data_master_read & ~onchip_memory2_1_s1_waits_for_read;

  //shift register p1 cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register = {cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register, cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in};

  //cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register <= 0;
      else 
        cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register <= p1_cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
    end


  //local readdatavalid cpu_2_data_master_read_data_valid_onchip_memory2_1_s1, which is an e_mux
  assign cpu_2_data_master_read_data_valid_onchip_memory2_1_s1 = cpu_2_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;

  assign cpu_2_instruction_master_requests_onchip_memory2_1_s1 = (({cpu_2_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h4000) & (cpu_2_instruction_master_read)) & cpu_2_instruction_master_read;
  assign cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1 = cpu_2_instruction_master_requests_onchip_memory2_1_s1 & ~((cpu_2_instruction_master_read & ((1 < cpu_2_instruction_master_latency_counter) | (|cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in = cpu_2_instruction_master_granted_onchip_memory2_1_s1 & cpu_2_instruction_master_read & ~onchip_memory2_1_s1_waits_for_read;

  //shift register p1 cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register = {cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register, cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in};

  //cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register <= 0;
      else 
        cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register <= p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
    end


  //local readdatavalid cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1, which is an e_mux
  assign cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1 = cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;

  assign cpu_3_data_master_requests_onchip_memory2_1_s1 = ({cpu_3_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h4000) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_onchip_memory2_1_s1 = cpu_3_data_master_requests_onchip_memory2_1_s1 & ~((cpu_3_data_master_read & ((1 < cpu_3_data_master_latency_counter) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in = cpu_3_data_master_granted_onchip_memory2_1_s1 & cpu_3_data_master_read & ~onchip_memory2_1_s1_waits_for_read;

  //shift register p1 cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register = {cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register, cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register_in};

  //cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register <= 0;
      else 
        cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register <= p1_cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;
    end


  //local readdatavalid cpu_3_data_master_read_data_valid_onchip_memory2_1_s1, which is an e_mux
  assign cpu_3_data_master_read_data_valid_onchip_memory2_1_s1 = cpu_3_data_master_read_data_valid_onchip_memory2_1_s1_shift_register;

  assign cpu_3_instruction_master_requests_onchip_memory2_1_s1 = (({cpu_3_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h4000) & (cpu_3_instruction_master_read)) & cpu_3_instruction_master_read;
  assign cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1 = cpu_3_instruction_master_requests_onchip_memory2_1_s1 & ~((cpu_3_instruction_master_read & ((1 < cpu_3_instruction_master_latency_counter) | (|cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in = cpu_3_instruction_master_granted_onchip_memory2_1_s1 & cpu_3_instruction_master_read & ~onchip_memory2_1_s1_waits_for_read;

  //shift register p1 cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register = {cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register, cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register_in};

  //cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register <= 0;
      else 
        cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register <= p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;
    end


  //local readdatavalid cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1, which is an e_mux
  assign cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1 = cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1_shift_register;

  //allow new arb cycle for onchip_memory2_1/s1, which is an e_assign
  assign onchip_memory2_1_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_1_instruction_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_2_instruction_master_arbiterlock & ~cpu_3_data_master_arbiterlock & ~cpu_3_instruction_master_arbiterlock;

  //cpu_3/instruction_master assignment into master qualified-requests vector for onchip_memory2_1/s1, which is an e_assign
  assign onchip_memory2_1_s1_master_qreq_vector[0] = cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1;

  //cpu_3/instruction_master grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_3_instruction_master_granted_onchip_memory2_1_s1 = onchip_memory2_1_s1_grant_vector[0];

  //cpu_3/instruction_master saved-grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_3_instruction_master_saved_grant_onchip_memory2_1_s1 = onchip_memory2_1_s1_arb_winner[0] && cpu_3_instruction_master_requests_onchip_memory2_1_s1;

  //cpu_3/data_master assignment into master qualified-requests vector for onchip_memory2_1/s1, which is an e_assign
  assign onchip_memory2_1_s1_master_qreq_vector[1] = cpu_3_data_master_qualified_request_onchip_memory2_1_s1;

  //cpu_3/data_master grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_3_data_master_granted_onchip_memory2_1_s1 = onchip_memory2_1_s1_grant_vector[1];

  //cpu_3/data_master saved-grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_3_data_master_saved_grant_onchip_memory2_1_s1 = onchip_memory2_1_s1_arb_winner[1] && cpu_3_data_master_requests_onchip_memory2_1_s1;

  //cpu_2/instruction_master assignment into master qualified-requests vector for onchip_memory2_1/s1, which is an e_assign
  assign onchip_memory2_1_s1_master_qreq_vector[2] = cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1;

  //cpu_2/instruction_master grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_2_instruction_master_granted_onchip_memory2_1_s1 = onchip_memory2_1_s1_grant_vector[2];

  //cpu_2/instruction_master saved-grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_2_instruction_master_saved_grant_onchip_memory2_1_s1 = onchip_memory2_1_s1_arb_winner[2] && cpu_2_instruction_master_requests_onchip_memory2_1_s1;

  //cpu_2/data_master assignment into master qualified-requests vector for onchip_memory2_1/s1, which is an e_assign
  assign onchip_memory2_1_s1_master_qreq_vector[3] = cpu_2_data_master_qualified_request_onchip_memory2_1_s1;

  //cpu_2/data_master grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_2_data_master_granted_onchip_memory2_1_s1 = onchip_memory2_1_s1_grant_vector[3];

  //cpu_2/data_master saved-grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_2_data_master_saved_grant_onchip_memory2_1_s1 = onchip_memory2_1_s1_arb_winner[3] && cpu_2_data_master_requests_onchip_memory2_1_s1;

  //cpu_1/instruction_master assignment into master qualified-requests vector for onchip_memory2_1/s1, which is an e_assign
  assign onchip_memory2_1_s1_master_qreq_vector[4] = cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1;

  //cpu_1/instruction_master grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_1_instruction_master_granted_onchip_memory2_1_s1 = onchip_memory2_1_s1_grant_vector[4];

  //cpu_1/instruction_master saved-grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_1_instruction_master_saved_grant_onchip_memory2_1_s1 = onchip_memory2_1_s1_arb_winner[4] && cpu_1_instruction_master_requests_onchip_memory2_1_s1;

  //cpu_1/data_master assignment into master qualified-requests vector for onchip_memory2_1/s1, which is an e_assign
  assign onchip_memory2_1_s1_master_qreq_vector[5] = cpu_1_data_master_qualified_request_onchip_memory2_1_s1;

  //cpu_1/data_master grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_1_data_master_granted_onchip_memory2_1_s1 = onchip_memory2_1_s1_grant_vector[5];

  //cpu_1/data_master saved-grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_1_data_master_saved_grant_onchip_memory2_1_s1 = onchip_memory2_1_s1_arb_winner[5] && cpu_1_data_master_requests_onchip_memory2_1_s1;

  //cpu_0/instruction_master assignment into master qualified-requests vector for onchip_memory2_1/s1, which is an e_assign
  assign onchip_memory2_1_s1_master_qreq_vector[6] = cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1;

  //cpu_0/instruction_master grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_0_instruction_master_granted_onchip_memory2_1_s1 = onchip_memory2_1_s1_grant_vector[6];

  //cpu_0/instruction_master saved-grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_onchip_memory2_1_s1 = onchip_memory2_1_s1_arb_winner[6] && cpu_0_instruction_master_requests_onchip_memory2_1_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for onchip_memory2_1/s1, which is an e_assign
  assign onchip_memory2_1_s1_master_qreq_vector[7] = cpu_0_data_master_qualified_request_onchip_memory2_1_s1;

  //cpu_0/data_master grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_0_data_master_granted_onchip_memory2_1_s1 = onchip_memory2_1_s1_grant_vector[7];

  //cpu_0/data_master saved-grant onchip_memory2_1/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_onchip_memory2_1_s1 = onchip_memory2_1_s1_arb_winner[7] && cpu_0_data_master_requests_onchip_memory2_1_s1;

  //onchip_memory2_1/s1 chosen-master double-vector, which is an e_assign
  assign onchip_memory2_1_s1_chosen_master_double_vector = {onchip_memory2_1_s1_master_qreq_vector, onchip_memory2_1_s1_master_qreq_vector} & ({~onchip_memory2_1_s1_master_qreq_vector, ~onchip_memory2_1_s1_master_qreq_vector} + onchip_memory2_1_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign onchip_memory2_1_s1_arb_winner = (onchip_memory2_1_s1_allow_new_arb_cycle & | onchip_memory2_1_s1_grant_vector) ? onchip_memory2_1_s1_grant_vector : onchip_memory2_1_s1_saved_chosen_master_vector;

  //saved onchip_memory2_1_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_1_s1_saved_chosen_master_vector <= 0;
      else if (onchip_memory2_1_s1_allow_new_arb_cycle)
          onchip_memory2_1_s1_saved_chosen_master_vector <= |onchip_memory2_1_s1_grant_vector ? onchip_memory2_1_s1_grant_vector : onchip_memory2_1_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign onchip_memory2_1_s1_grant_vector = {(onchip_memory2_1_s1_chosen_master_double_vector[7] | onchip_memory2_1_s1_chosen_master_double_vector[15]),
    (onchip_memory2_1_s1_chosen_master_double_vector[6] | onchip_memory2_1_s1_chosen_master_double_vector[14]),
    (onchip_memory2_1_s1_chosen_master_double_vector[5] | onchip_memory2_1_s1_chosen_master_double_vector[13]),
    (onchip_memory2_1_s1_chosen_master_double_vector[4] | onchip_memory2_1_s1_chosen_master_double_vector[12]),
    (onchip_memory2_1_s1_chosen_master_double_vector[3] | onchip_memory2_1_s1_chosen_master_double_vector[11]),
    (onchip_memory2_1_s1_chosen_master_double_vector[2] | onchip_memory2_1_s1_chosen_master_double_vector[10]),
    (onchip_memory2_1_s1_chosen_master_double_vector[1] | onchip_memory2_1_s1_chosen_master_double_vector[9]),
    (onchip_memory2_1_s1_chosen_master_double_vector[0] | onchip_memory2_1_s1_chosen_master_double_vector[8])};

  //onchip_memory2_1/s1 chosen master rotated left, which is an e_assign
  assign onchip_memory2_1_s1_chosen_master_rot_left = (onchip_memory2_1_s1_arb_winner << 1) ? (onchip_memory2_1_s1_arb_winner << 1) : 1;

  //onchip_memory2_1/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_1_s1_arb_addend <= 1;
      else if (|onchip_memory2_1_s1_grant_vector)
          onchip_memory2_1_s1_arb_addend <= onchip_memory2_1_s1_end_xfer? onchip_memory2_1_s1_chosen_master_rot_left : onchip_memory2_1_s1_grant_vector;
    end


  //~onchip_memory2_1_s1_reset assignment, which is an e_assign
  assign onchip_memory2_1_s1_reset = ~reset_n;

  assign onchip_memory2_1_s1_chipselect = cpu_0_data_master_granted_onchip_memory2_1_s1 | cpu_0_instruction_master_granted_onchip_memory2_1_s1 | cpu_1_data_master_granted_onchip_memory2_1_s1 | cpu_1_instruction_master_granted_onchip_memory2_1_s1 | cpu_2_data_master_granted_onchip_memory2_1_s1 | cpu_2_instruction_master_granted_onchip_memory2_1_s1 | cpu_3_data_master_granted_onchip_memory2_1_s1 | cpu_3_instruction_master_granted_onchip_memory2_1_s1;
  //onchip_memory2_1_s1_firsttransfer first transaction, which is an e_assign
  assign onchip_memory2_1_s1_firsttransfer = onchip_memory2_1_s1_begins_xfer ? onchip_memory2_1_s1_unreg_firsttransfer : onchip_memory2_1_s1_reg_firsttransfer;

  //onchip_memory2_1_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign onchip_memory2_1_s1_unreg_firsttransfer = ~(onchip_memory2_1_s1_slavearbiterlockenable & onchip_memory2_1_s1_any_continuerequest);

  //onchip_memory2_1_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_1_s1_reg_firsttransfer <= 1'b1;
      else if (onchip_memory2_1_s1_begins_xfer)
          onchip_memory2_1_s1_reg_firsttransfer <= onchip_memory2_1_s1_unreg_firsttransfer;
    end


  //onchip_memory2_1_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign onchip_memory2_1_s1_beginbursttransfer_internal = onchip_memory2_1_s1_begins_xfer;

  //onchip_memory2_1_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign onchip_memory2_1_s1_arbitration_holdoff_internal = onchip_memory2_1_s1_begins_xfer & onchip_memory2_1_s1_firsttransfer;

  //onchip_memory2_1_s1_write assignment, which is an e_mux
  assign onchip_memory2_1_s1_write = (cpu_0_data_master_granted_onchip_memory2_1_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_onchip_memory2_1_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_onchip_memory2_1_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_onchip_memory2_1_s1 & cpu_3_data_master_write);

  assign shifted_address_to_onchip_memory2_1_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //onchip_memory2_1_s1_address mux, which is an e_mux
  assign onchip_memory2_1_s1_address = (cpu_0_data_master_granted_onchip_memory2_1_s1)? (shifted_address_to_onchip_memory2_1_s1_from_cpu_0_data_master >> 2) :
    (cpu_0_instruction_master_granted_onchip_memory2_1_s1)? (shifted_address_to_onchip_memory2_1_s1_from_cpu_0_instruction_master >> 2) :
    (cpu_1_data_master_granted_onchip_memory2_1_s1)? (shifted_address_to_onchip_memory2_1_s1_from_cpu_1_data_master >> 2) :
    (cpu_1_instruction_master_granted_onchip_memory2_1_s1)? (shifted_address_to_onchip_memory2_1_s1_from_cpu_1_instruction_master >> 2) :
    (cpu_2_data_master_granted_onchip_memory2_1_s1)? (shifted_address_to_onchip_memory2_1_s1_from_cpu_2_data_master >> 2) :
    (cpu_2_instruction_master_granted_onchip_memory2_1_s1)? (shifted_address_to_onchip_memory2_1_s1_from_cpu_2_instruction_master >> 2) :
    (cpu_3_data_master_granted_onchip_memory2_1_s1)? (shifted_address_to_onchip_memory2_1_s1_from_cpu_3_data_master >> 2) :
    (shifted_address_to_onchip_memory2_1_s1_from_cpu_3_instruction_master >> 2);

  assign shifted_address_to_onchip_memory2_1_s1_from_cpu_0_instruction_master = cpu_0_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_1_s1_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_1_s1_from_cpu_1_instruction_master = cpu_1_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_1_s1_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_1_s1_from_cpu_2_instruction_master = cpu_2_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_1_s1_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_1_s1_from_cpu_3_instruction_master = cpu_3_instruction_master_address_to_slave;
  //d1_onchip_memory2_1_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_onchip_memory2_1_s1_end_xfer <= 1;
      else 
        d1_onchip_memory2_1_s1_end_xfer <= onchip_memory2_1_s1_end_xfer;
    end


  //onchip_memory2_1_s1_waits_for_read in a cycle, which is an e_mux
  assign onchip_memory2_1_s1_waits_for_read = onchip_memory2_1_s1_in_a_read_cycle & 0;

  //onchip_memory2_1_s1_in_a_read_cycle assignment, which is an e_assign
  assign onchip_memory2_1_s1_in_a_read_cycle = (cpu_0_data_master_granted_onchip_memory2_1_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_onchip_memory2_1_s1 & cpu_0_instruction_master_read) | (cpu_1_data_master_granted_onchip_memory2_1_s1 & cpu_1_data_master_read) | (cpu_1_instruction_master_granted_onchip_memory2_1_s1 & cpu_1_instruction_master_read) | (cpu_2_data_master_granted_onchip_memory2_1_s1 & cpu_2_data_master_read) | (cpu_2_instruction_master_granted_onchip_memory2_1_s1 & cpu_2_instruction_master_read) | (cpu_3_data_master_granted_onchip_memory2_1_s1 & cpu_3_data_master_read) | (cpu_3_instruction_master_granted_onchip_memory2_1_s1 & cpu_3_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = onchip_memory2_1_s1_in_a_read_cycle;

  //onchip_memory2_1_s1_waits_for_write in a cycle, which is an e_mux
  assign onchip_memory2_1_s1_waits_for_write = onchip_memory2_1_s1_in_a_write_cycle & 0;

  //onchip_memory2_1_s1_in_a_write_cycle assignment, which is an e_assign
  assign onchip_memory2_1_s1_in_a_write_cycle = (cpu_0_data_master_granted_onchip_memory2_1_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_onchip_memory2_1_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_onchip_memory2_1_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_onchip_memory2_1_s1 & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = onchip_memory2_1_s1_in_a_write_cycle;

  assign wait_for_onchip_memory2_1_s1_counter = 0;
  //onchip_memory2_1_s1_byteenable byte enable port mux, which is an e_mux
  assign onchip_memory2_1_s1_byteenable = (cpu_0_data_master_granted_onchip_memory2_1_s1)? cpu_0_data_master_byteenable :
    (cpu_1_data_master_granted_onchip_memory2_1_s1)? cpu_1_data_master_byteenable :
    (cpu_2_data_master_granted_onchip_memory2_1_s1)? cpu_2_data_master_byteenable :
    (cpu_3_data_master_granted_onchip_memory2_1_s1)? cpu_3_data_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //onchip_memory2_1/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_onchip_memory2_1_s1 + cpu_0_instruction_master_granted_onchip_memory2_1_s1 + cpu_1_data_master_granted_onchip_memory2_1_s1 + cpu_1_instruction_master_granted_onchip_memory2_1_s1 + cpu_2_data_master_granted_onchip_memory2_1_s1 + cpu_2_instruction_master_granted_onchip_memory2_1_s1 + cpu_3_data_master_granted_onchip_memory2_1_s1 + cpu_3_instruction_master_granted_onchip_memory2_1_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_onchip_memory2_1_s1 + cpu_0_instruction_master_saved_grant_onchip_memory2_1_s1 + cpu_1_data_master_saved_grant_onchip_memory2_1_s1 + cpu_1_instruction_master_saved_grant_onchip_memory2_1_s1 + cpu_2_data_master_saved_grant_onchip_memory2_1_s1 + cpu_2_instruction_master_saved_grant_onchip_memory2_1_s1 + cpu_3_data_master_saved_grant_onchip_memory2_1_s1 + cpu_3_instruction_master_saved_grant_onchip_memory2_1_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module onchip_memory2_2_s1_arbitrator (
                                        // inputs:
                                         clk,
                                         cpu_0_data_master_address_to_slave,
                                         cpu_0_data_master_byteenable,
                                         cpu_0_data_master_latency_counter,
                                         cpu_0_data_master_read,
                                         cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_0_data_master_write,
                                         cpu_0_data_master_writedata,
                                         cpu_0_instruction_master_address_to_slave,
                                         cpu_0_instruction_master_latency_counter,
                                         cpu_0_instruction_master_read,
                                         cpu_1_data_master_address_to_slave,
                                         cpu_1_data_master_byteenable,
                                         cpu_1_data_master_latency_counter,
                                         cpu_1_data_master_read,
                                         cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_1_data_master_write,
                                         cpu_1_data_master_writedata,
                                         cpu_1_instruction_master_address_to_slave,
                                         cpu_1_instruction_master_latency_counter,
                                         cpu_1_instruction_master_read,
                                         cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_2_data_master_address_to_slave,
                                         cpu_2_data_master_byteenable,
                                         cpu_2_data_master_latency_counter,
                                         cpu_2_data_master_read,
                                         cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_2_data_master_write,
                                         cpu_2_data_master_writedata,
                                         cpu_2_instruction_master_address_to_slave,
                                         cpu_2_instruction_master_latency_counter,
                                         cpu_2_instruction_master_read,
                                         cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_3_data_master_address_to_slave,
                                         cpu_3_data_master_byteenable,
                                         cpu_3_data_master_latency_counter,
                                         cpu_3_data_master_read,
                                         cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_3_data_master_write,
                                         cpu_3_data_master_writedata,
                                         cpu_3_instruction_master_address_to_slave,
                                         cpu_3_instruction_master_latency_counter,
                                         cpu_3_instruction_master_read,
                                         cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         onchip_memory2_2_s1_readdata,
                                         reset_n,

                                        // outputs:
                                         cpu_0_data_master_granted_onchip_memory2_2_s1,
                                         cpu_0_data_master_qualified_request_onchip_memory2_2_s1,
                                         cpu_0_data_master_read_data_valid_onchip_memory2_2_s1,
                                         cpu_0_data_master_requests_onchip_memory2_2_s1,
                                         cpu_0_instruction_master_granted_onchip_memory2_2_s1,
                                         cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1,
                                         cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1,
                                         cpu_0_instruction_master_requests_onchip_memory2_2_s1,
                                         cpu_1_data_master_granted_onchip_memory2_2_s1,
                                         cpu_1_data_master_qualified_request_onchip_memory2_2_s1,
                                         cpu_1_data_master_read_data_valid_onchip_memory2_2_s1,
                                         cpu_1_data_master_requests_onchip_memory2_2_s1,
                                         cpu_1_instruction_master_granted_onchip_memory2_2_s1,
                                         cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1,
                                         cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1,
                                         cpu_1_instruction_master_requests_onchip_memory2_2_s1,
                                         cpu_2_data_master_granted_onchip_memory2_2_s1,
                                         cpu_2_data_master_qualified_request_onchip_memory2_2_s1,
                                         cpu_2_data_master_read_data_valid_onchip_memory2_2_s1,
                                         cpu_2_data_master_requests_onchip_memory2_2_s1,
                                         cpu_2_instruction_master_granted_onchip_memory2_2_s1,
                                         cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1,
                                         cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1,
                                         cpu_2_instruction_master_requests_onchip_memory2_2_s1,
                                         cpu_3_data_master_granted_onchip_memory2_2_s1,
                                         cpu_3_data_master_qualified_request_onchip_memory2_2_s1,
                                         cpu_3_data_master_read_data_valid_onchip_memory2_2_s1,
                                         cpu_3_data_master_requests_onchip_memory2_2_s1,
                                         cpu_3_instruction_master_granted_onchip_memory2_2_s1,
                                         cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1,
                                         cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1,
                                         cpu_3_instruction_master_requests_onchip_memory2_2_s1,
                                         d1_onchip_memory2_2_s1_end_xfer,
                                         onchip_memory2_2_s1_address,
                                         onchip_memory2_2_s1_byteenable,
                                         onchip_memory2_2_s1_chipselect,
                                         onchip_memory2_2_s1_clken,
                                         onchip_memory2_2_s1_readdata_from_sa,
                                         onchip_memory2_2_s1_reset,
                                         onchip_memory2_2_s1_write,
                                         onchip_memory2_2_s1_writedata
                                      )
;

  output           cpu_0_data_master_granted_onchip_memory2_2_s1;
  output           cpu_0_data_master_qualified_request_onchip_memory2_2_s1;
  output           cpu_0_data_master_read_data_valid_onchip_memory2_2_s1;
  output           cpu_0_data_master_requests_onchip_memory2_2_s1;
  output           cpu_0_instruction_master_granted_onchip_memory2_2_s1;
  output           cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1;
  output           cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1;
  output           cpu_0_instruction_master_requests_onchip_memory2_2_s1;
  output           cpu_1_data_master_granted_onchip_memory2_2_s1;
  output           cpu_1_data_master_qualified_request_onchip_memory2_2_s1;
  output           cpu_1_data_master_read_data_valid_onchip_memory2_2_s1;
  output           cpu_1_data_master_requests_onchip_memory2_2_s1;
  output           cpu_1_instruction_master_granted_onchip_memory2_2_s1;
  output           cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1;
  output           cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1;
  output           cpu_1_instruction_master_requests_onchip_memory2_2_s1;
  output           cpu_2_data_master_granted_onchip_memory2_2_s1;
  output           cpu_2_data_master_qualified_request_onchip_memory2_2_s1;
  output           cpu_2_data_master_read_data_valid_onchip_memory2_2_s1;
  output           cpu_2_data_master_requests_onchip_memory2_2_s1;
  output           cpu_2_instruction_master_granted_onchip_memory2_2_s1;
  output           cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1;
  output           cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1;
  output           cpu_2_instruction_master_requests_onchip_memory2_2_s1;
  output           cpu_3_data_master_granted_onchip_memory2_2_s1;
  output           cpu_3_data_master_qualified_request_onchip_memory2_2_s1;
  output           cpu_3_data_master_read_data_valid_onchip_memory2_2_s1;
  output           cpu_3_data_master_requests_onchip_memory2_2_s1;
  output           cpu_3_instruction_master_granted_onchip_memory2_2_s1;
  output           cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1;
  output           cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1;
  output           cpu_3_instruction_master_requests_onchip_memory2_2_s1;
  output           d1_onchip_memory2_2_s1_end_xfer;
  output  [  6: 0] onchip_memory2_2_s1_address;
  output  [  3: 0] onchip_memory2_2_s1_byteenable;
  output           onchip_memory2_2_s1_chipselect;
  output           onchip_memory2_2_s1_clken;
  output  [ 31: 0] onchip_memory2_2_s1_readdata_from_sa;
  output           onchip_memory2_2_s1_reset;
  output           onchip_memory2_2_s1_write;
  output  [ 31: 0] onchip_memory2_2_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input            cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input   [  3: 0] cpu_1_data_master_byteenable;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_1_instruction_master_address_to_slave;
  input            cpu_1_instruction_master_latency_counter;
  input            cpu_1_instruction_master_read;
  input            cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input   [  3: 0] cpu_2_data_master_byteenable;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_2_instruction_master_address_to_slave;
  input            cpu_2_instruction_master_latency_counter;
  input            cpu_2_instruction_master_read;
  input            cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input   [  3: 0] cpu_3_data_master_byteenable;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 24: 0] cpu_3_instruction_master_address_to_slave;
  input            cpu_3_instruction_master_latency_counter;
  input            cpu_3_instruction_master_read;
  input            cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 31: 0] onchip_memory2_2_s1_readdata;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_onchip_memory2_2_s1;
  wire             cpu_0_data_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_2_s1;
  reg              cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in;
  wire             cpu_0_data_master_requests_onchip_memory2_2_s1;
  wire             cpu_0_data_master_saved_grant_onchip_memory2_2_s1;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_onchip_memory2_2_s1;
  wire             cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1;
  reg              cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in;
  wire             cpu_0_instruction_master_requests_onchip_memory2_2_s1;
  wire             cpu_0_instruction_master_saved_grant_onchip_memory2_2_s1;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_onchip_memory2_2_s1;
  wire             cpu_1_data_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_2_s1;
  reg              cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in;
  wire             cpu_1_data_master_requests_onchip_memory2_2_s1;
  wire             cpu_1_data_master_saved_grant_onchip_memory2_2_s1;
  wire             cpu_1_instruction_master_arbiterlock;
  wire             cpu_1_instruction_master_arbiterlock2;
  wire             cpu_1_instruction_master_continuerequest;
  wire             cpu_1_instruction_master_granted_onchip_memory2_2_s1;
  wire             cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1;
  reg              cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in;
  wire             cpu_1_instruction_master_requests_onchip_memory2_2_s1;
  wire             cpu_1_instruction_master_saved_grant_onchip_memory2_2_s1;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_onchip_memory2_2_s1;
  wire             cpu_2_data_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_2_s1;
  reg              cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in;
  wire             cpu_2_data_master_requests_onchip_memory2_2_s1;
  wire             cpu_2_data_master_saved_grant_onchip_memory2_2_s1;
  wire             cpu_2_instruction_master_arbiterlock;
  wire             cpu_2_instruction_master_arbiterlock2;
  wire             cpu_2_instruction_master_continuerequest;
  wire             cpu_2_instruction_master_granted_onchip_memory2_2_s1;
  wire             cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1;
  reg              cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in;
  wire             cpu_2_instruction_master_requests_onchip_memory2_2_s1;
  wire             cpu_2_instruction_master_saved_grant_onchip_memory2_2_s1;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_onchip_memory2_2_s1;
  wire             cpu_3_data_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_2_s1;
  reg              cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in;
  wire             cpu_3_data_master_requests_onchip_memory2_2_s1;
  wire             cpu_3_data_master_saved_grant_onchip_memory2_2_s1;
  wire             cpu_3_instruction_master_arbiterlock;
  wire             cpu_3_instruction_master_arbiterlock2;
  wire             cpu_3_instruction_master_continuerequest;
  wire             cpu_3_instruction_master_granted_onchip_memory2_2_s1;
  wire             cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1;
  reg              cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in;
  wire             cpu_3_instruction_master_requests_onchip_memory2_2_s1;
  wire             cpu_3_instruction_master_saved_grant_onchip_memory2_2_s1;
  reg              d1_onchip_memory2_2_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_onchip_memory2_2_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_2_s1;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_2_s1;
  reg              last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_2_s1;
  reg              last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_2_s1;
  reg              last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_2_s1;
  reg              last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_2_s1;
  reg              last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_2_s1;
  reg              last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_2_s1;
  wire    [  6: 0] onchip_memory2_2_s1_address;
  wire             onchip_memory2_2_s1_allgrants;
  wire             onchip_memory2_2_s1_allow_new_arb_cycle;
  wire             onchip_memory2_2_s1_any_bursting_master_saved_grant;
  wire             onchip_memory2_2_s1_any_continuerequest;
  reg     [  7: 0] onchip_memory2_2_s1_arb_addend;
  wire             onchip_memory2_2_s1_arb_counter_enable;
  reg     [  2: 0] onchip_memory2_2_s1_arb_share_counter;
  wire    [  2: 0] onchip_memory2_2_s1_arb_share_counter_next_value;
  wire    [  2: 0] onchip_memory2_2_s1_arb_share_set_values;
  wire    [  7: 0] onchip_memory2_2_s1_arb_winner;
  wire             onchip_memory2_2_s1_arbitration_holdoff_internal;
  wire             onchip_memory2_2_s1_beginbursttransfer_internal;
  wire             onchip_memory2_2_s1_begins_xfer;
  wire    [  3: 0] onchip_memory2_2_s1_byteenable;
  wire             onchip_memory2_2_s1_chipselect;
  wire    [ 15: 0] onchip_memory2_2_s1_chosen_master_double_vector;
  wire    [  7: 0] onchip_memory2_2_s1_chosen_master_rot_left;
  wire             onchip_memory2_2_s1_clken;
  wire             onchip_memory2_2_s1_end_xfer;
  wire             onchip_memory2_2_s1_firsttransfer;
  wire    [  7: 0] onchip_memory2_2_s1_grant_vector;
  wire             onchip_memory2_2_s1_in_a_read_cycle;
  wire             onchip_memory2_2_s1_in_a_write_cycle;
  wire    [  7: 0] onchip_memory2_2_s1_master_qreq_vector;
  wire             onchip_memory2_2_s1_non_bursting_master_requests;
  wire    [ 31: 0] onchip_memory2_2_s1_readdata_from_sa;
  reg              onchip_memory2_2_s1_reg_firsttransfer;
  wire             onchip_memory2_2_s1_reset;
  reg     [  7: 0] onchip_memory2_2_s1_saved_chosen_master_vector;
  reg              onchip_memory2_2_s1_slavearbiterlockenable;
  wire             onchip_memory2_2_s1_slavearbiterlockenable2;
  wire             onchip_memory2_2_s1_unreg_firsttransfer;
  wire             onchip_memory2_2_s1_waits_for_read;
  wire             onchip_memory2_2_s1_waits_for_write;
  wire             onchip_memory2_2_s1_write;
  wire    [ 31: 0] onchip_memory2_2_s1_writedata;
  wire             p1_cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             p1_cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             p1_cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             p1_cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire             p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_2_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_2_s1_from_cpu_0_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_2_s1_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_2_s1_from_cpu_1_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_2_s1_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_2_s1_from_cpu_2_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_2_s1_from_cpu_3_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_2_s1_from_cpu_3_instruction_master;
  wire             wait_for_onchip_memory2_2_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~onchip_memory2_2_s1_end_xfer;
    end


  assign onchip_memory2_2_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_onchip_memory2_2_s1 | cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1 | cpu_1_data_master_qualified_request_onchip_memory2_2_s1 | cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1 | cpu_2_data_master_qualified_request_onchip_memory2_2_s1 | cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1 | cpu_3_data_master_qualified_request_onchip_memory2_2_s1 | cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1));
  //assign onchip_memory2_2_s1_readdata_from_sa = onchip_memory2_2_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign onchip_memory2_2_s1_readdata_from_sa = onchip_memory2_2_s1_readdata;

  assign cpu_0_data_master_requests_onchip_memory2_2_s1 = ({cpu_0_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h6000) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //onchip_memory2_2_s1_arb_share_counter set values, which is an e_mux
  assign onchip_memory2_2_s1_arb_share_set_values = 1;

  //onchip_memory2_2_s1_non_bursting_master_requests mux, which is an e_mux
  assign onchip_memory2_2_s1_non_bursting_master_requests = cpu_0_data_master_requests_onchip_memory2_2_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_1_data_master_requests_onchip_memory2_2_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_2_data_master_requests_onchip_memory2_2_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_3_data_master_requests_onchip_memory2_2_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_0_data_master_requests_onchip_memory2_2_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_1_data_master_requests_onchip_memory2_2_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_2_data_master_requests_onchip_memory2_2_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_3_data_master_requests_onchip_memory2_2_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_0_data_master_requests_onchip_memory2_2_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_1_data_master_requests_onchip_memory2_2_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_2_data_master_requests_onchip_memory2_2_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_3_data_master_requests_onchip_memory2_2_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_0_data_master_requests_onchip_memory2_2_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_1_data_master_requests_onchip_memory2_2_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_2_data_master_requests_onchip_memory2_2_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_3_data_master_requests_onchip_memory2_2_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_0_data_master_requests_onchip_memory2_2_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_1_data_master_requests_onchip_memory2_2_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_2_data_master_requests_onchip_memory2_2_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_3_data_master_requests_onchip_memory2_2_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_0_data_master_requests_onchip_memory2_2_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_1_data_master_requests_onchip_memory2_2_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_2_data_master_requests_onchip_memory2_2_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_3_data_master_requests_onchip_memory2_2_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_0_data_master_requests_onchip_memory2_2_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_1_data_master_requests_onchip_memory2_2_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_2_data_master_requests_onchip_memory2_2_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_3_data_master_requests_onchip_memory2_2_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_0_data_master_requests_onchip_memory2_2_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_1_data_master_requests_onchip_memory2_2_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_2_data_master_requests_onchip_memory2_2_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_2_s1 |
    cpu_3_data_master_requests_onchip_memory2_2_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_2_s1;

  //onchip_memory2_2_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign onchip_memory2_2_s1_any_bursting_master_saved_grant = 0;

  //onchip_memory2_2_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign onchip_memory2_2_s1_arb_share_counter_next_value = onchip_memory2_2_s1_firsttransfer ? (onchip_memory2_2_s1_arb_share_set_values - 1) : |onchip_memory2_2_s1_arb_share_counter ? (onchip_memory2_2_s1_arb_share_counter - 1) : 0;

  //onchip_memory2_2_s1_allgrants all slave grants, which is an e_mux
  assign onchip_memory2_2_s1_allgrants = (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector) |
    (|onchip_memory2_2_s1_grant_vector);

  //onchip_memory2_2_s1_end_xfer assignment, which is an e_assign
  assign onchip_memory2_2_s1_end_xfer = ~(onchip_memory2_2_s1_waits_for_read | onchip_memory2_2_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_onchip_memory2_2_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_onchip_memory2_2_s1 = onchip_memory2_2_s1_end_xfer & (~onchip_memory2_2_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //onchip_memory2_2_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign onchip_memory2_2_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_onchip_memory2_2_s1 & onchip_memory2_2_s1_allgrants) | (end_xfer_arb_share_counter_term_onchip_memory2_2_s1 & ~onchip_memory2_2_s1_non_bursting_master_requests);

  //onchip_memory2_2_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_2_s1_arb_share_counter <= 0;
      else if (onchip_memory2_2_s1_arb_counter_enable)
          onchip_memory2_2_s1_arb_share_counter <= onchip_memory2_2_s1_arb_share_counter_next_value;
    end


  //onchip_memory2_2_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_2_s1_slavearbiterlockenable <= 0;
      else if ((|onchip_memory2_2_s1_master_qreq_vector & end_xfer_arb_share_counter_term_onchip_memory2_2_s1) | (end_xfer_arb_share_counter_term_onchip_memory2_2_s1 & ~onchip_memory2_2_s1_non_bursting_master_requests))
          onchip_memory2_2_s1_slavearbiterlockenable <= |onchip_memory2_2_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master onchip_memory2_2/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = onchip_memory2_2_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //onchip_memory2_2_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign onchip_memory2_2_s1_slavearbiterlockenable2 = |onchip_memory2_2_s1_arb_share_counter_next_value;

  //cpu_0/data_master onchip_memory2_2/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = onchip_memory2_2_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master onchip_memory2_2/s1 arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = onchip_memory2_2_s1_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master onchip_memory2_2/s1 arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = onchip_memory2_2_s1_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted onchip_memory2_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_2_s1 <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_2_s1 <= cpu_0_instruction_master_saved_grant_onchip_memory2_2_s1 ? 1 : (onchip_memory2_2_s1_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_onchip_memory2_2_s1) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_2_s1;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_0_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_0_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_0_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_0_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_0_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_0_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_0_instruction_master_requests_onchip_memory2_2_s1);

  //onchip_memory2_2_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign onchip_memory2_2_s1_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest;

  //cpu_1/data_master onchip_memory2_2/s1 arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = onchip_memory2_2_s1_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master onchip_memory2_2/s1 arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = onchip_memory2_2_s1_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted onchip_memory2_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_2_s1 <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_2_s1 <= cpu_1_data_master_saved_grant_onchip_memory2_2_s1 ? 1 : (onchip_memory2_2_s1_arbitration_holdoff_internal | ~cpu_1_data_master_requests_onchip_memory2_2_s1) ? 0 : last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_2_s1;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_2_s1 & cpu_1_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_2_s1 & cpu_1_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_2_s1 & cpu_1_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_2_s1 & cpu_1_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_2_s1 & cpu_1_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_2_s1 & cpu_1_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_2_s1 & cpu_1_data_master_requests_onchip_memory2_2_s1);

  //cpu_1/instruction_master onchip_memory2_2/s1 arbiterlock, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock = onchip_memory2_2_s1_slavearbiterlockenable & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master onchip_memory2_2/s1 arbiterlock2, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock2 = onchip_memory2_2_s1_slavearbiterlockenable2 & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master granted onchip_memory2_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_2_s1 <= 0;
      else 
        last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_2_s1 <= cpu_1_instruction_master_saved_grant_onchip_memory2_2_s1 ? 1 : (onchip_memory2_2_s1_arbitration_holdoff_internal | ~cpu_1_instruction_master_requests_onchip_memory2_2_s1) ? 0 : last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_2_s1;
    end


  //cpu_1_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_1_instruction_master_continuerequest = (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_1_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_1_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_1_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_1_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_1_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_1_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_1_instruction_master_requests_onchip_memory2_2_s1);

  //cpu_2/data_master onchip_memory2_2/s1 arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = onchip_memory2_2_s1_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master onchip_memory2_2/s1 arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = onchip_memory2_2_s1_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted onchip_memory2_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_2_s1 <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_2_s1 <= cpu_2_data_master_saved_grant_onchip_memory2_2_s1 ? 1 : (onchip_memory2_2_s1_arbitration_holdoff_internal | ~cpu_2_data_master_requests_onchip_memory2_2_s1) ? 0 : last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_2_s1;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_2_s1 & cpu_2_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_2_s1 & cpu_2_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_2_s1 & cpu_2_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_2_s1 & cpu_2_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_2_s1 & cpu_2_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_2_s1 & cpu_2_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_2_s1 & cpu_2_data_master_requests_onchip_memory2_2_s1);

  //cpu_2/instruction_master onchip_memory2_2/s1 arbiterlock, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock = onchip_memory2_2_s1_slavearbiterlockenable & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master onchip_memory2_2/s1 arbiterlock2, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock2 = onchip_memory2_2_s1_slavearbiterlockenable2 & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master granted onchip_memory2_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_2_s1 <= 0;
      else 
        last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_2_s1 <= cpu_2_instruction_master_saved_grant_onchip_memory2_2_s1 ? 1 : (onchip_memory2_2_s1_arbitration_holdoff_internal | ~cpu_2_instruction_master_requests_onchip_memory2_2_s1) ? 0 : last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_2_s1;
    end


  //cpu_2_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_2_instruction_master_continuerequest = (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_2_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_2_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_2_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_2_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_2_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_2_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_2_instruction_master_requests_onchip_memory2_2_s1);

  //cpu_3/data_master onchip_memory2_2/s1 arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = onchip_memory2_2_s1_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master onchip_memory2_2/s1 arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = onchip_memory2_2_s1_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted onchip_memory2_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_2_s1 <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_2_s1 <= cpu_3_data_master_saved_grant_onchip_memory2_2_s1 ? 1 : (onchip_memory2_2_s1_arbitration_holdoff_internal | ~cpu_3_data_master_requests_onchip_memory2_2_s1) ? 0 : last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_2_s1;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_2_s1 & cpu_3_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_2_s1 & cpu_3_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_2_s1 & cpu_3_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_2_s1 & cpu_3_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_2_s1 & cpu_3_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_2_s1 & cpu_3_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_2_s1 & cpu_3_data_master_requests_onchip_memory2_2_s1);

  //cpu_3/instruction_master onchip_memory2_2/s1 arbiterlock, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock = onchip_memory2_2_s1_slavearbiterlockenable & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master onchip_memory2_2/s1 arbiterlock2, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock2 = onchip_memory2_2_s1_slavearbiterlockenable2 & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master granted onchip_memory2_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_2_s1 <= 0;
      else 
        last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_2_s1 <= cpu_3_instruction_master_saved_grant_onchip_memory2_2_s1 ? 1 : (onchip_memory2_2_s1_arbitration_holdoff_internal | ~cpu_3_instruction_master_requests_onchip_memory2_2_s1) ? 0 : last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_2_s1;
    end


  //cpu_3_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_3_instruction_master_continuerequest = (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_3_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_3_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_3_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_3_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_3_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_3_instruction_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_2_s1 & cpu_3_instruction_master_requests_onchip_memory2_2_s1);

  assign cpu_0_data_master_qualified_request_onchip_memory2_2_s1 = cpu_0_data_master_requests_onchip_memory2_2_s1 & ~((cpu_0_data_master_read & ((1 < cpu_0_data_master_latency_counter) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in = cpu_0_data_master_granted_onchip_memory2_2_s1 & cpu_0_data_master_read & ~onchip_memory2_2_s1_waits_for_read;

  //shift register p1 cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register = {cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register, cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in};

  //cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register <= 0;
      else 
        cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register <= p1_cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
    end


  //local readdatavalid cpu_0_data_master_read_data_valid_onchip_memory2_2_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_onchip_memory2_2_s1 = cpu_0_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;

  //onchip_memory2_2_s1_writedata mux, which is an e_mux
  assign onchip_memory2_2_s1_writedata = (cpu_0_data_master_granted_onchip_memory2_2_s1)? cpu_0_data_master_writedata :
    (cpu_1_data_master_granted_onchip_memory2_2_s1)? cpu_1_data_master_writedata :
    (cpu_2_data_master_granted_onchip_memory2_2_s1)? cpu_2_data_master_writedata :
    cpu_3_data_master_writedata;

  //mux onchip_memory2_2_s1_clken, which is an e_mux
  assign onchip_memory2_2_s1_clken = 1'b1;

  assign cpu_0_instruction_master_requests_onchip_memory2_2_s1 = (({cpu_0_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h6000) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted onchip_memory2_2/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_2_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_2_s1 <= cpu_0_data_master_saved_grant_onchip_memory2_2_s1 ? 1 : (onchip_memory2_2_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_onchip_memory2_2_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_2_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_2_s1 & cpu_0_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_2_s1 & cpu_0_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_2_s1 & cpu_0_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_2_s1 & cpu_0_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_2_s1 & cpu_0_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_2_s1 & cpu_0_data_master_requests_onchip_memory2_2_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_2_s1 & cpu_0_data_master_requests_onchip_memory2_2_s1);

  assign cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1 = cpu_0_instruction_master_requests_onchip_memory2_2_s1 & ~((cpu_0_instruction_master_read & ((1 < cpu_0_instruction_master_latency_counter))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in = cpu_0_instruction_master_granted_onchip_memory2_2_s1 & cpu_0_instruction_master_read & ~onchip_memory2_2_s1_waits_for_read;

  //shift register p1 cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register = {cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register, cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in};

  //cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register <= 0;
      else 
        cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register <= p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
    end


  //local readdatavalid cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1 = cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;

  assign cpu_1_data_master_requests_onchip_memory2_2_s1 = ({cpu_1_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h6000) & (cpu_1_data_master_read | cpu_1_data_master_write);
  assign cpu_1_data_master_qualified_request_onchip_memory2_2_s1 = cpu_1_data_master_requests_onchip_memory2_2_s1 & ~((cpu_1_data_master_read & ((1 < cpu_1_data_master_latency_counter) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in = cpu_1_data_master_granted_onchip_memory2_2_s1 & cpu_1_data_master_read & ~onchip_memory2_2_s1_waits_for_read;

  //shift register p1 cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register = {cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register, cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in};

  //cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register <= 0;
      else 
        cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register <= p1_cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
    end


  //local readdatavalid cpu_1_data_master_read_data_valid_onchip_memory2_2_s1, which is an e_mux
  assign cpu_1_data_master_read_data_valid_onchip_memory2_2_s1 = cpu_1_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;

  assign cpu_1_instruction_master_requests_onchip_memory2_2_s1 = (({cpu_1_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h6000) & (cpu_1_instruction_master_read)) & cpu_1_instruction_master_read;
  assign cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1 = cpu_1_instruction_master_requests_onchip_memory2_2_s1 & ~((cpu_1_instruction_master_read & ((1 < cpu_1_instruction_master_latency_counter) | (|cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in = cpu_1_instruction_master_granted_onchip_memory2_2_s1 & cpu_1_instruction_master_read & ~onchip_memory2_2_s1_waits_for_read;

  //shift register p1 cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register = {cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register, cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in};

  //cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register <= 0;
      else 
        cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register <= p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
    end


  //local readdatavalid cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1, which is an e_mux
  assign cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1 = cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;

  assign cpu_2_data_master_requests_onchip_memory2_2_s1 = ({cpu_2_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h6000) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_onchip_memory2_2_s1 = cpu_2_data_master_requests_onchip_memory2_2_s1 & ~((cpu_2_data_master_read & ((1 < cpu_2_data_master_latency_counter) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in = cpu_2_data_master_granted_onchip_memory2_2_s1 & cpu_2_data_master_read & ~onchip_memory2_2_s1_waits_for_read;

  //shift register p1 cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register = {cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register, cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in};

  //cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register <= 0;
      else 
        cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register <= p1_cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
    end


  //local readdatavalid cpu_2_data_master_read_data_valid_onchip_memory2_2_s1, which is an e_mux
  assign cpu_2_data_master_read_data_valid_onchip_memory2_2_s1 = cpu_2_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;

  assign cpu_2_instruction_master_requests_onchip_memory2_2_s1 = (({cpu_2_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h6000) & (cpu_2_instruction_master_read)) & cpu_2_instruction_master_read;
  assign cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1 = cpu_2_instruction_master_requests_onchip_memory2_2_s1 & ~((cpu_2_instruction_master_read & ((1 < cpu_2_instruction_master_latency_counter) | (|cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in = cpu_2_instruction_master_granted_onchip_memory2_2_s1 & cpu_2_instruction_master_read & ~onchip_memory2_2_s1_waits_for_read;

  //shift register p1 cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register = {cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register, cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in};

  //cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register <= 0;
      else 
        cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register <= p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
    end


  //local readdatavalid cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1, which is an e_mux
  assign cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1 = cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;

  assign cpu_3_data_master_requests_onchip_memory2_2_s1 = ({cpu_3_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h6000) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_onchip_memory2_2_s1 = cpu_3_data_master_requests_onchip_memory2_2_s1 & ~((cpu_3_data_master_read & ((1 < cpu_3_data_master_latency_counter) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in = cpu_3_data_master_granted_onchip_memory2_2_s1 & cpu_3_data_master_read & ~onchip_memory2_2_s1_waits_for_read;

  //shift register p1 cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register = {cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register, cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register_in};

  //cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register <= 0;
      else 
        cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register <= p1_cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;
    end


  //local readdatavalid cpu_3_data_master_read_data_valid_onchip_memory2_2_s1, which is an e_mux
  assign cpu_3_data_master_read_data_valid_onchip_memory2_2_s1 = cpu_3_data_master_read_data_valid_onchip_memory2_2_s1_shift_register;

  assign cpu_3_instruction_master_requests_onchip_memory2_2_s1 = (({cpu_3_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h6000) & (cpu_3_instruction_master_read)) & cpu_3_instruction_master_read;
  assign cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1 = cpu_3_instruction_master_requests_onchip_memory2_2_s1 & ~((cpu_3_instruction_master_read & ((1 < cpu_3_instruction_master_latency_counter) | (|cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in = cpu_3_instruction_master_granted_onchip_memory2_2_s1 & cpu_3_instruction_master_read & ~onchip_memory2_2_s1_waits_for_read;

  //shift register p1 cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register = {cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register, cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register_in};

  //cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register <= 0;
      else 
        cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register <= p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;
    end


  //local readdatavalid cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1, which is an e_mux
  assign cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1 = cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1_shift_register;

  //allow new arb cycle for onchip_memory2_2/s1, which is an e_assign
  assign onchip_memory2_2_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_1_instruction_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_2_instruction_master_arbiterlock & ~cpu_3_data_master_arbiterlock & ~cpu_3_instruction_master_arbiterlock;

  //cpu_3/instruction_master assignment into master qualified-requests vector for onchip_memory2_2/s1, which is an e_assign
  assign onchip_memory2_2_s1_master_qreq_vector[0] = cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1;

  //cpu_3/instruction_master grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_3_instruction_master_granted_onchip_memory2_2_s1 = onchip_memory2_2_s1_grant_vector[0];

  //cpu_3/instruction_master saved-grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_3_instruction_master_saved_grant_onchip_memory2_2_s1 = onchip_memory2_2_s1_arb_winner[0] && cpu_3_instruction_master_requests_onchip_memory2_2_s1;

  //cpu_3/data_master assignment into master qualified-requests vector for onchip_memory2_2/s1, which is an e_assign
  assign onchip_memory2_2_s1_master_qreq_vector[1] = cpu_3_data_master_qualified_request_onchip_memory2_2_s1;

  //cpu_3/data_master grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_3_data_master_granted_onchip_memory2_2_s1 = onchip_memory2_2_s1_grant_vector[1];

  //cpu_3/data_master saved-grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_3_data_master_saved_grant_onchip_memory2_2_s1 = onchip_memory2_2_s1_arb_winner[1] && cpu_3_data_master_requests_onchip_memory2_2_s1;

  //cpu_2/instruction_master assignment into master qualified-requests vector for onchip_memory2_2/s1, which is an e_assign
  assign onchip_memory2_2_s1_master_qreq_vector[2] = cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1;

  //cpu_2/instruction_master grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_2_instruction_master_granted_onchip_memory2_2_s1 = onchip_memory2_2_s1_grant_vector[2];

  //cpu_2/instruction_master saved-grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_2_instruction_master_saved_grant_onchip_memory2_2_s1 = onchip_memory2_2_s1_arb_winner[2] && cpu_2_instruction_master_requests_onchip_memory2_2_s1;

  //cpu_2/data_master assignment into master qualified-requests vector for onchip_memory2_2/s1, which is an e_assign
  assign onchip_memory2_2_s1_master_qreq_vector[3] = cpu_2_data_master_qualified_request_onchip_memory2_2_s1;

  //cpu_2/data_master grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_2_data_master_granted_onchip_memory2_2_s1 = onchip_memory2_2_s1_grant_vector[3];

  //cpu_2/data_master saved-grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_2_data_master_saved_grant_onchip_memory2_2_s1 = onchip_memory2_2_s1_arb_winner[3] && cpu_2_data_master_requests_onchip_memory2_2_s1;

  //cpu_1/instruction_master assignment into master qualified-requests vector for onchip_memory2_2/s1, which is an e_assign
  assign onchip_memory2_2_s1_master_qreq_vector[4] = cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1;

  //cpu_1/instruction_master grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_1_instruction_master_granted_onchip_memory2_2_s1 = onchip_memory2_2_s1_grant_vector[4];

  //cpu_1/instruction_master saved-grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_1_instruction_master_saved_grant_onchip_memory2_2_s1 = onchip_memory2_2_s1_arb_winner[4] && cpu_1_instruction_master_requests_onchip_memory2_2_s1;

  //cpu_1/data_master assignment into master qualified-requests vector for onchip_memory2_2/s1, which is an e_assign
  assign onchip_memory2_2_s1_master_qreq_vector[5] = cpu_1_data_master_qualified_request_onchip_memory2_2_s1;

  //cpu_1/data_master grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_1_data_master_granted_onchip_memory2_2_s1 = onchip_memory2_2_s1_grant_vector[5];

  //cpu_1/data_master saved-grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_1_data_master_saved_grant_onchip_memory2_2_s1 = onchip_memory2_2_s1_arb_winner[5] && cpu_1_data_master_requests_onchip_memory2_2_s1;

  //cpu_0/instruction_master assignment into master qualified-requests vector for onchip_memory2_2/s1, which is an e_assign
  assign onchip_memory2_2_s1_master_qreq_vector[6] = cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1;

  //cpu_0/instruction_master grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_0_instruction_master_granted_onchip_memory2_2_s1 = onchip_memory2_2_s1_grant_vector[6];

  //cpu_0/instruction_master saved-grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_onchip_memory2_2_s1 = onchip_memory2_2_s1_arb_winner[6] && cpu_0_instruction_master_requests_onchip_memory2_2_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for onchip_memory2_2/s1, which is an e_assign
  assign onchip_memory2_2_s1_master_qreq_vector[7] = cpu_0_data_master_qualified_request_onchip_memory2_2_s1;

  //cpu_0/data_master grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_0_data_master_granted_onchip_memory2_2_s1 = onchip_memory2_2_s1_grant_vector[7];

  //cpu_0/data_master saved-grant onchip_memory2_2/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_onchip_memory2_2_s1 = onchip_memory2_2_s1_arb_winner[7] && cpu_0_data_master_requests_onchip_memory2_2_s1;

  //onchip_memory2_2/s1 chosen-master double-vector, which is an e_assign
  assign onchip_memory2_2_s1_chosen_master_double_vector = {onchip_memory2_2_s1_master_qreq_vector, onchip_memory2_2_s1_master_qreq_vector} & ({~onchip_memory2_2_s1_master_qreq_vector, ~onchip_memory2_2_s1_master_qreq_vector} + onchip_memory2_2_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign onchip_memory2_2_s1_arb_winner = (onchip_memory2_2_s1_allow_new_arb_cycle & | onchip_memory2_2_s1_grant_vector) ? onchip_memory2_2_s1_grant_vector : onchip_memory2_2_s1_saved_chosen_master_vector;

  //saved onchip_memory2_2_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_2_s1_saved_chosen_master_vector <= 0;
      else if (onchip_memory2_2_s1_allow_new_arb_cycle)
          onchip_memory2_2_s1_saved_chosen_master_vector <= |onchip_memory2_2_s1_grant_vector ? onchip_memory2_2_s1_grant_vector : onchip_memory2_2_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign onchip_memory2_2_s1_grant_vector = {(onchip_memory2_2_s1_chosen_master_double_vector[7] | onchip_memory2_2_s1_chosen_master_double_vector[15]),
    (onchip_memory2_2_s1_chosen_master_double_vector[6] | onchip_memory2_2_s1_chosen_master_double_vector[14]),
    (onchip_memory2_2_s1_chosen_master_double_vector[5] | onchip_memory2_2_s1_chosen_master_double_vector[13]),
    (onchip_memory2_2_s1_chosen_master_double_vector[4] | onchip_memory2_2_s1_chosen_master_double_vector[12]),
    (onchip_memory2_2_s1_chosen_master_double_vector[3] | onchip_memory2_2_s1_chosen_master_double_vector[11]),
    (onchip_memory2_2_s1_chosen_master_double_vector[2] | onchip_memory2_2_s1_chosen_master_double_vector[10]),
    (onchip_memory2_2_s1_chosen_master_double_vector[1] | onchip_memory2_2_s1_chosen_master_double_vector[9]),
    (onchip_memory2_2_s1_chosen_master_double_vector[0] | onchip_memory2_2_s1_chosen_master_double_vector[8])};

  //onchip_memory2_2/s1 chosen master rotated left, which is an e_assign
  assign onchip_memory2_2_s1_chosen_master_rot_left = (onchip_memory2_2_s1_arb_winner << 1) ? (onchip_memory2_2_s1_arb_winner << 1) : 1;

  //onchip_memory2_2/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_2_s1_arb_addend <= 1;
      else if (|onchip_memory2_2_s1_grant_vector)
          onchip_memory2_2_s1_arb_addend <= onchip_memory2_2_s1_end_xfer? onchip_memory2_2_s1_chosen_master_rot_left : onchip_memory2_2_s1_grant_vector;
    end


  //~onchip_memory2_2_s1_reset assignment, which is an e_assign
  assign onchip_memory2_2_s1_reset = ~reset_n;

  assign onchip_memory2_2_s1_chipselect = cpu_0_data_master_granted_onchip_memory2_2_s1 | cpu_0_instruction_master_granted_onchip_memory2_2_s1 | cpu_1_data_master_granted_onchip_memory2_2_s1 | cpu_1_instruction_master_granted_onchip_memory2_2_s1 | cpu_2_data_master_granted_onchip_memory2_2_s1 | cpu_2_instruction_master_granted_onchip_memory2_2_s1 | cpu_3_data_master_granted_onchip_memory2_2_s1 | cpu_3_instruction_master_granted_onchip_memory2_2_s1;
  //onchip_memory2_2_s1_firsttransfer first transaction, which is an e_assign
  assign onchip_memory2_2_s1_firsttransfer = onchip_memory2_2_s1_begins_xfer ? onchip_memory2_2_s1_unreg_firsttransfer : onchip_memory2_2_s1_reg_firsttransfer;

  //onchip_memory2_2_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign onchip_memory2_2_s1_unreg_firsttransfer = ~(onchip_memory2_2_s1_slavearbiterlockenable & onchip_memory2_2_s1_any_continuerequest);

  //onchip_memory2_2_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_2_s1_reg_firsttransfer <= 1'b1;
      else if (onchip_memory2_2_s1_begins_xfer)
          onchip_memory2_2_s1_reg_firsttransfer <= onchip_memory2_2_s1_unreg_firsttransfer;
    end


  //onchip_memory2_2_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign onchip_memory2_2_s1_beginbursttransfer_internal = onchip_memory2_2_s1_begins_xfer;

  //onchip_memory2_2_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign onchip_memory2_2_s1_arbitration_holdoff_internal = onchip_memory2_2_s1_begins_xfer & onchip_memory2_2_s1_firsttransfer;

  //onchip_memory2_2_s1_write assignment, which is an e_mux
  assign onchip_memory2_2_s1_write = (cpu_0_data_master_granted_onchip_memory2_2_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_onchip_memory2_2_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_onchip_memory2_2_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_onchip_memory2_2_s1 & cpu_3_data_master_write);

  assign shifted_address_to_onchip_memory2_2_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //onchip_memory2_2_s1_address mux, which is an e_mux
  assign onchip_memory2_2_s1_address = (cpu_0_data_master_granted_onchip_memory2_2_s1)? (shifted_address_to_onchip_memory2_2_s1_from_cpu_0_data_master >> 2) :
    (cpu_0_instruction_master_granted_onchip_memory2_2_s1)? (shifted_address_to_onchip_memory2_2_s1_from_cpu_0_instruction_master >> 2) :
    (cpu_1_data_master_granted_onchip_memory2_2_s1)? (shifted_address_to_onchip_memory2_2_s1_from_cpu_1_data_master >> 2) :
    (cpu_1_instruction_master_granted_onchip_memory2_2_s1)? (shifted_address_to_onchip_memory2_2_s1_from_cpu_1_instruction_master >> 2) :
    (cpu_2_data_master_granted_onchip_memory2_2_s1)? (shifted_address_to_onchip_memory2_2_s1_from_cpu_2_data_master >> 2) :
    (cpu_2_instruction_master_granted_onchip_memory2_2_s1)? (shifted_address_to_onchip_memory2_2_s1_from_cpu_2_instruction_master >> 2) :
    (cpu_3_data_master_granted_onchip_memory2_2_s1)? (shifted_address_to_onchip_memory2_2_s1_from_cpu_3_data_master >> 2) :
    (shifted_address_to_onchip_memory2_2_s1_from_cpu_3_instruction_master >> 2);

  assign shifted_address_to_onchip_memory2_2_s1_from_cpu_0_instruction_master = cpu_0_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_2_s1_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_2_s1_from_cpu_1_instruction_master = cpu_1_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_2_s1_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_2_s1_from_cpu_2_instruction_master = cpu_2_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_2_s1_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_2_s1_from_cpu_3_instruction_master = cpu_3_instruction_master_address_to_slave;
  //d1_onchip_memory2_2_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_onchip_memory2_2_s1_end_xfer <= 1;
      else 
        d1_onchip_memory2_2_s1_end_xfer <= onchip_memory2_2_s1_end_xfer;
    end


  //onchip_memory2_2_s1_waits_for_read in a cycle, which is an e_mux
  assign onchip_memory2_2_s1_waits_for_read = onchip_memory2_2_s1_in_a_read_cycle & 0;

  //onchip_memory2_2_s1_in_a_read_cycle assignment, which is an e_assign
  assign onchip_memory2_2_s1_in_a_read_cycle = (cpu_0_data_master_granted_onchip_memory2_2_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_onchip_memory2_2_s1 & cpu_0_instruction_master_read) | (cpu_1_data_master_granted_onchip_memory2_2_s1 & cpu_1_data_master_read) | (cpu_1_instruction_master_granted_onchip_memory2_2_s1 & cpu_1_instruction_master_read) | (cpu_2_data_master_granted_onchip_memory2_2_s1 & cpu_2_data_master_read) | (cpu_2_instruction_master_granted_onchip_memory2_2_s1 & cpu_2_instruction_master_read) | (cpu_3_data_master_granted_onchip_memory2_2_s1 & cpu_3_data_master_read) | (cpu_3_instruction_master_granted_onchip_memory2_2_s1 & cpu_3_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = onchip_memory2_2_s1_in_a_read_cycle;

  //onchip_memory2_2_s1_waits_for_write in a cycle, which is an e_mux
  assign onchip_memory2_2_s1_waits_for_write = onchip_memory2_2_s1_in_a_write_cycle & 0;

  //onchip_memory2_2_s1_in_a_write_cycle assignment, which is an e_assign
  assign onchip_memory2_2_s1_in_a_write_cycle = (cpu_0_data_master_granted_onchip_memory2_2_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_onchip_memory2_2_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_onchip_memory2_2_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_onchip_memory2_2_s1 & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = onchip_memory2_2_s1_in_a_write_cycle;

  assign wait_for_onchip_memory2_2_s1_counter = 0;
  //onchip_memory2_2_s1_byteenable byte enable port mux, which is an e_mux
  assign onchip_memory2_2_s1_byteenable = (cpu_0_data_master_granted_onchip_memory2_2_s1)? cpu_0_data_master_byteenable :
    (cpu_1_data_master_granted_onchip_memory2_2_s1)? cpu_1_data_master_byteenable :
    (cpu_2_data_master_granted_onchip_memory2_2_s1)? cpu_2_data_master_byteenable :
    (cpu_3_data_master_granted_onchip_memory2_2_s1)? cpu_3_data_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //onchip_memory2_2/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_onchip_memory2_2_s1 + cpu_0_instruction_master_granted_onchip_memory2_2_s1 + cpu_1_data_master_granted_onchip_memory2_2_s1 + cpu_1_instruction_master_granted_onchip_memory2_2_s1 + cpu_2_data_master_granted_onchip_memory2_2_s1 + cpu_2_instruction_master_granted_onchip_memory2_2_s1 + cpu_3_data_master_granted_onchip_memory2_2_s1 + cpu_3_instruction_master_granted_onchip_memory2_2_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_onchip_memory2_2_s1 + cpu_0_instruction_master_saved_grant_onchip_memory2_2_s1 + cpu_1_data_master_saved_grant_onchip_memory2_2_s1 + cpu_1_instruction_master_saved_grant_onchip_memory2_2_s1 + cpu_2_data_master_saved_grant_onchip_memory2_2_s1 + cpu_2_instruction_master_saved_grant_onchip_memory2_2_s1 + cpu_3_data_master_saved_grant_onchip_memory2_2_s1 + cpu_3_instruction_master_saved_grant_onchip_memory2_2_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module onchip_memory2_3_s1_arbitrator (
                                        // inputs:
                                         clk,
                                         cpu_0_data_master_address_to_slave,
                                         cpu_0_data_master_byteenable,
                                         cpu_0_data_master_latency_counter,
                                         cpu_0_data_master_read,
                                         cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_0_data_master_write,
                                         cpu_0_data_master_writedata,
                                         cpu_0_instruction_master_address_to_slave,
                                         cpu_0_instruction_master_latency_counter,
                                         cpu_0_instruction_master_read,
                                         cpu_1_data_master_address_to_slave,
                                         cpu_1_data_master_byteenable,
                                         cpu_1_data_master_latency_counter,
                                         cpu_1_data_master_read,
                                         cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_1_data_master_write,
                                         cpu_1_data_master_writedata,
                                         cpu_1_instruction_master_address_to_slave,
                                         cpu_1_instruction_master_latency_counter,
                                         cpu_1_instruction_master_read,
                                         cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_2_data_master_address_to_slave,
                                         cpu_2_data_master_byteenable,
                                         cpu_2_data_master_latency_counter,
                                         cpu_2_data_master_read,
                                         cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_2_data_master_write,
                                         cpu_2_data_master_writedata,
                                         cpu_2_instruction_master_address_to_slave,
                                         cpu_2_instruction_master_latency_counter,
                                         cpu_2_instruction_master_read,
                                         cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_3_data_master_address_to_slave,
                                         cpu_3_data_master_byteenable,
                                         cpu_3_data_master_latency_counter,
                                         cpu_3_data_master_read,
                                         cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_3_data_master_write,
                                         cpu_3_data_master_writedata,
                                         cpu_3_instruction_master_address_to_slave,
                                         cpu_3_instruction_master_latency_counter,
                                         cpu_3_instruction_master_read,
                                         cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         onchip_memory2_3_s1_readdata,
                                         reset_n,

                                        // outputs:
                                         cpu_0_data_master_granted_onchip_memory2_3_s1,
                                         cpu_0_data_master_qualified_request_onchip_memory2_3_s1,
                                         cpu_0_data_master_read_data_valid_onchip_memory2_3_s1,
                                         cpu_0_data_master_requests_onchip_memory2_3_s1,
                                         cpu_0_instruction_master_granted_onchip_memory2_3_s1,
                                         cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1,
                                         cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1,
                                         cpu_0_instruction_master_requests_onchip_memory2_3_s1,
                                         cpu_1_data_master_granted_onchip_memory2_3_s1,
                                         cpu_1_data_master_qualified_request_onchip_memory2_3_s1,
                                         cpu_1_data_master_read_data_valid_onchip_memory2_3_s1,
                                         cpu_1_data_master_requests_onchip_memory2_3_s1,
                                         cpu_1_instruction_master_granted_onchip_memory2_3_s1,
                                         cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1,
                                         cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1,
                                         cpu_1_instruction_master_requests_onchip_memory2_3_s1,
                                         cpu_2_data_master_granted_onchip_memory2_3_s1,
                                         cpu_2_data_master_qualified_request_onchip_memory2_3_s1,
                                         cpu_2_data_master_read_data_valid_onchip_memory2_3_s1,
                                         cpu_2_data_master_requests_onchip_memory2_3_s1,
                                         cpu_2_instruction_master_granted_onchip_memory2_3_s1,
                                         cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1,
                                         cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1,
                                         cpu_2_instruction_master_requests_onchip_memory2_3_s1,
                                         cpu_3_data_master_granted_onchip_memory2_3_s1,
                                         cpu_3_data_master_qualified_request_onchip_memory2_3_s1,
                                         cpu_3_data_master_read_data_valid_onchip_memory2_3_s1,
                                         cpu_3_data_master_requests_onchip_memory2_3_s1,
                                         cpu_3_instruction_master_granted_onchip_memory2_3_s1,
                                         cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1,
                                         cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1,
                                         cpu_3_instruction_master_requests_onchip_memory2_3_s1,
                                         d1_onchip_memory2_3_s1_end_xfer,
                                         onchip_memory2_3_s1_address,
                                         onchip_memory2_3_s1_byteenable,
                                         onchip_memory2_3_s1_chipselect,
                                         onchip_memory2_3_s1_clken,
                                         onchip_memory2_3_s1_readdata_from_sa,
                                         onchip_memory2_3_s1_reset,
                                         onchip_memory2_3_s1_write,
                                         onchip_memory2_3_s1_writedata
                                      )
;

  output           cpu_0_data_master_granted_onchip_memory2_3_s1;
  output           cpu_0_data_master_qualified_request_onchip_memory2_3_s1;
  output           cpu_0_data_master_read_data_valid_onchip_memory2_3_s1;
  output           cpu_0_data_master_requests_onchip_memory2_3_s1;
  output           cpu_0_instruction_master_granted_onchip_memory2_3_s1;
  output           cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1;
  output           cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1;
  output           cpu_0_instruction_master_requests_onchip_memory2_3_s1;
  output           cpu_1_data_master_granted_onchip_memory2_3_s1;
  output           cpu_1_data_master_qualified_request_onchip_memory2_3_s1;
  output           cpu_1_data_master_read_data_valid_onchip_memory2_3_s1;
  output           cpu_1_data_master_requests_onchip_memory2_3_s1;
  output           cpu_1_instruction_master_granted_onchip_memory2_3_s1;
  output           cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1;
  output           cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1;
  output           cpu_1_instruction_master_requests_onchip_memory2_3_s1;
  output           cpu_2_data_master_granted_onchip_memory2_3_s1;
  output           cpu_2_data_master_qualified_request_onchip_memory2_3_s1;
  output           cpu_2_data_master_read_data_valid_onchip_memory2_3_s1;
  output           cpu_2_data_master_requests_onchip_memory2_3_s1;
  output           cpu_2_instruction_master_granted_onchip_memory2_3_s1;
  output           cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1;
  output           cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1;
  output           cpu_2_instruction_master_requests_onchip_memory2_3_s1;
  output           cpu_3_data_master_granted_onchip_memory2_3_s1;
  output           cpu_3_data_master_qualified_request_onchip_memory2_3_s1;
  output           cpu_3_data_master_read_data_valid_onchip_memory2_3_s1;
  output           cpu_3_data_master_requests_onchip_memory2_3_s1;
  output           cpu_3_instruction_master_granted_onchip_memory2_3_s1;
  output           cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1;
  output           cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1;
  output           cpu_3_instruction_master_requests_onchip_memory2_3_s1;
  output           d1_onchip_memory2_3_s1_end_xfer;
  output  [  6: 0] onchip_memory2_3_s1_address;
  output  [  3: 0] onchip_memory2_3_s1_byteenable;
  output           onchip_memory2_3_s1_chipselect;
  output           onchip_memory2_3_s1_clken;
  output  [ 31: 0] onchip_memory2_3_s1_readdata_from_sa;
  output           onchip_memory2_3_s1_reset;
  output           onchip_memory2_3_s1_write;
  output  [ 31: 0] onchip_memory2_3_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input            cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input   [  3: 0] cpu_1_data_master_byteenable;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_1_instruction_master_address_to_slave;
  input            cpu_1_instruction_master_latency_counter;
  input            cpu_1_instruction_master_read;
  input            cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input   [  3: 0] cpu_2_data_master_byteenable;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_2_instruction_master_address_to_slave;
  input            cpu_2_instruction_master_latency_counter;
  input            cpu_2_instruction_master_read;
  input            cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input   [  3: 0] cpu_3_data_master_byteenable;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 24: 0] cpu_3_instruction_master_address_to_slave;
  input            cpu_3_instruction_master_latency_counter;
  input            cpu_3_instruction_master_read;
  input            cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input   [ 31: 0] onchip_memory2_3_s1_readdata;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_onchip_memory2_3_s1;
  wire             cpu_0_data_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_3_s1;
  reg              cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in;
  wire             cpu_0_data_master_requests_onchip_memory2_3_s1;
  wire             cpu_0_data_master_saved_grant_onchip_memory2_3_s1;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_onchip_memory2_3_s1;
  wire             cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1;
  reg              cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in;
  wire             cpu_0_instruction_master_requests_onchip_memory2_3_s1;
  wire             cpu_0_instruction_master_saved_grant_onchip_memory2_3_s1;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_onchip_memory2_3_s1;
  wire             cpu_1_data_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_3_s1;
  reg              cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in;
  wire             cpu_1_data_master_requests_onchip_memory2_3_s1;
  wire             cpu_1_data_master_saved_grant_onchip_memory2_3_s1;
  wire             cpu_1_instruction_master_arbiterlock;
  wire             cpu_1_instruction_master_arbiterlock2;
  wire             cpu_1_instruction_master_continuerequest;
  wire             cpu_1_instruction_master_granted_onchip_memory2_3_s1;
  wire             cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1;
  reg              cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in;
  wire             cpu_1_instruction_master_requests_onchip_memory2_3_s1;
  wire             cpu_1_instruction_master_saved_grant_onchip_memory2_3_s1;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_onchip_memory2_3_s1;
  wire             cpu_2_data_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_3_s1;
  reg              cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in;
  wire             cpu_2_data_master_requests_onchip_memory2_3_s1;
  wire             cpu_2_data_master_saved_grant_onchip_memory2_3_s1;
  wire             cpu_2_instruction_master_arbiterlock;
  wire             cpu_2_instruction_master_arbiterlock2;
  wire             cpu_2_instruction_master_continuerequest;
  wire             cpu_2_instruction_master_granted_onchip_memory2_3_s1;
  wire             cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1;
  reg              cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in;
  wire             cpu_2_instruction_master_requests_onchip_memory2_3_s1;
  wire             cpu_2_instruction_master_saved_grant_onchip_memory2_3_s1;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_onchip_memory2_3_s1;
  wire             cpu_3_data_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_3_s1;
  reg              cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in;
  wire             cpu_3_data_master_requests_onchip_memory2_3_s1;
  wire             cpu_3_data_master_saved_grant_onchip_memory2_3_s1;
  wire             cpu_3_instruction_master_arbiterlock;
  wire             cpu_3_instruction_master_arbiterlock2;
  wire             cpu_3_instruction_master_continuerequest;
  wire             cpu_3_instruction_master_granted_onchip_memory2_3_s1;
  wire             cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1;
  reg              cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in;
  wire             cpu_3_instruction_master_requests_onchip_memory2_3_s1;
  wire             cpu_3_instruction_master_saved_grant_onchip_memory2_3_s1;
  reg              d1_onchip_memory2_3_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_onchip_memory2_3_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_3_s1;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_3_s1;
  reg              last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_3_s1;
  reg              last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_3_s1;
  reg              last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_3_s1;
  reg              last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_3_s1;
  reg              last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_3_s1;
  reg              last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_3_s1;
  wire    [  6: 0] onchip_memory2_3_s1_address;
  wire             onchip_memory2_3_s1_allgrants;
  wire             onchip_memory2_3_s1_allow_new_arb_cycle;
  wire             onchip_memory2_3_s1_any_bursting_master_saved_grant;
  wire             onchip_memory2_3_s1_any_continuerequest;
  reg     [  7: 0] onchip_memory2_3_s1_arb_addend;
  wire             onchip_memory2_3_s1_arb_counter_enable;
  reg     [  2: 0] onchip_memory2_3_s1_arb_share_counter;
  wire    [  2: 0] onchip_memory2_3_s1_arb_share_counter_next_value;
  wire    [  2: 0] onchip_memory2_3_s1_arb_share_set_values;
  wire    [  7: 0] onchip_memory2_3_s1_arb_winner;
  wire             onchip_memory2_3_s1_arbitration_holdoff_internal;
  wire             onchip_memory2_3_s1_beginbursttransfer_internal;
  wire             onchip_memory2_3_s1_begins_xfer;
  wire    [  3: 0] onchip_memory2_3_s1_byteenable;
  wire             onchip_memory2_3_s1_chipselect;
  wire    [ 15: 0] onchip_memory2_3_s1_chosen_master_double_vector;
  wire    [  7: 0] onchip_memory2_3_s1_chosen_master_rot_left;
  wire             onchip_memory2_3_s1_clken;
  wire             onchip_memory2_3_s1_end_xfer;
  wire             onchip_memory2_3_s1_firsttransfer;
  wire    [  7: 0] onchip_memory2_3_s1_grant_vector;
  wire             onchip_memory2_3_s1_in_a_read_cycle;
  wire             onchip_memory2_3_s1_in_a_write_cycle;
  wire    [  7: 0] onchip_memory2_3_s1_master_qreq_vector;
  wire             onchip_memory2_3_s1_non_bursting_master_requests;
  wire    [ 31: 0] onchip_memory2_3_s1_readdata_from_sa;
  reg              onchip_memory2_3_s1_reg_firsttransfer;
  wire             onchip_memory2_3_s1_reset;
  reg     [  7: 0] onchip_memory2_3_s1_saved_chosen_master_vector;
  reg              onchip_memory2_3_s1_slavearbiterlockenable;
  wire             onchip_memory2_3_s1_slavearbiterlockenable2;
  wire             onchip_memory2_3_s1_unreg_firsttransfer;
  wire             onchip_memory2_3_s1_waits_for_read;
  wire             onchip_memory2_3_s1_waits_for_write;
  wire             onchip_memory2_3_s1_write;
  wire    [ 31: 0] onchip_memory2_3_s1_writedata;
  wire             p1_cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             p1_cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             p1_cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             p1_cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire             p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_3_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_3_s1_from_cpu_0_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_3_s1_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_3_s1_from_cpu_1_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_3_s1_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_3_s1_from_cpu_2_instruction_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_3_s1_from_cpu_3_data_master;
  wire    [ 24: 0] shifted_address_to_onchip_memory2_3_s1_from_cpu_3_instruction_master;
  wire             wait_for_onchip_memory2_3_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~onchip_memory2_3_s1_end_xfer;
    end


  assign onchip_memory2_3_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_onchip_memory2_3_s1 | cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1 | cpu_1_data_master_qualified_request_onchip_memory2_3_s1 | cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1 | cpu_2_data_master_qualified_request_onchip_memory2_3_s1 | cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1 | cpu_3_data_master_qualified_request_onchip_memory2_3_s1 | cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1));
  //assign onchip_memory2_3_s1_readdata_from_sa = onchip_memory2_3_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign onchip_memory2_3_s1_readdata_from_sa = onchip_memory2_3_s1_readdata;

  assign cpu_0_data_master_requests_onchip_memory2_3_s1 = ({cpu_0_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h7000) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //onchip_memory2_3_s1_arb_share_counter set values, which is an e_mux
  assign onchip_memory2_3_s1_arb_share_set_values = 1;

  //onchip_memory2_3_s1_non_bursting_master_requests mux, which is an e_mux
  assign onchip_memory2_3_s1_non_bursting_master_requests = cpu_0_data_master_requests_onchip_memory2_3_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_1_data_master_requests_onchip_memory2_3_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_2_data_master_requests_onchip_memory2_3_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_3_data_master_requests_onchip_memory2_3_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_0_data_master_requests_onchip_memory2_3_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_1_data_master_requests_onchip_memory2_3_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_2_data_master_requests_onchip_memory2_3_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_3_data_master_requests_onchip_memory2_3_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_0_data_master_requests_onchip_memory2_3_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_1_data_master_requests_onchip_memory2_3_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_2_data_master_requests_onchip_memory2_3_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_3_data_master_requests_onchip_memory2_3_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_0_data_master_requests_onchip_memory2_3_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_1_data_master_requests_onchip_memory2_3_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_2_data_master_requests_onchip_memory2_3_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_3_data_master_requests_onchip_memory2_3_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_0_data_master_requests_onchip_memory2_3_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_1_data_master_requests_onchip_memory2_3_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_2_data_master_requests_onchip_memory2_3_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_3_data_master_requests_onchip_memory2_3_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_0_data_master_requests_onchip_memory2_3_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_1_data_master_requests_onchip_memory2_3_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_2_data_master_requests_onchip_memory2_3_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_3_data_master_requests_onchip_memory2_3_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_0_data_master_requests_onchip_memory2_3_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_1_data_master_requests_onchip_memory2_3_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_2_data_master_requests_onchip_memory2_3_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_3_data_master_requests_onchip_memory2_3_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_0_data_master_requests_onchip_memory2_3_s1 |
    cpu_0_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_1_data_master_requests_onchip_memory2_3_s1 |
    cpu_1_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_2_data_master_requests_onchip_memory2_3_s1 |
    cpu_2_instruction_master_requests_onchip_memory2_3_s1 |
    cpu_3_data_master_requests_onchip_memory2_3_s1 |
    cpu_3_instruction_master_requests_onchip_memory2_3_s1;

  //onchip_memory2_3_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign onchip_memory2_3_s1_any_bursting_master_saved_grant = 0;

  //onchip_memory2_3_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign onchip_memory2_3_s1_arb_share_counter_next_value = onchip_memory2_3_s1_firsttransfer ? (onchip_memory2_3_s1_arb_share_set_values - 1) : |onchip_memory2_3_s1_arb_share_counter ? (onchip_memory2_3_s1_arb_share_counter - 1) : 0;

  //onchip_memory2_3_s1_allgrants all slave grants, which is an e_mux
  assign onchip_memory2_3_s1_allgrants = (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector) |
    (|onchip_memory2_3_s1_grant_vector);

  //onchip_memory2_3_s1_end_xfer assignment, which is an e_assign
  assign onchip_memory2_3_s1_end_xfer = ~(onchip_memory2_3_s1_waits_for_read | onchip_memory2_3_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_onchip_memory2_3_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_onchip_memory2_3_s1 = onchip_memory2_3_s1_end_xfer & (~onchip_memory2_3_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //onchip_memory2_3_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign onchip_memory2_3_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_onchip_memory2_3_s1 & onchip_memory2_3_s1_allgrants) | (end_xfer_arb_share_counter_term_onchip_memory2_3_s1 & ~onchip_memory2_3_s1_non_bursting_master_requests);

  //onchip_memory2_3_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_3_s1_arb_share_counter <= 0;
      else if (onchip_memory2_3_s1_arb_counter_enable)
          onchip_memory2_3_s1_arb_share_counter <= onchip_memory2_3_s1_arb_share_counter_next_value;
    end


  //onchip_memory2_3_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_3_s1_slavearbiterlockenable <= 0;
      else if ((|onchip_memory2_3_s1_master_qreq_vector & end_xfer_arb_share_counter_term_onchip_memory2_3_s1) | (end_xfer_arb_share_counter_term_onchip_memory2_3_s1 & ~onchip_memory2_3_s1_non_bursting_master_requests))
          onchip_memory2_3_s1_slavearbiterlockenable <= |onchip_memory2_3_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master onchip_memory2_3/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = onchip_memory2_3_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //onchip_memory2_3_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign onchip_memory2_3_s1_slavearbiterlockenable2 = |onchip_memory2_3_s1_arb_share_counter_next_value;

  //cpu_0/data_master onchip_memory2_3/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = onchip_memory2_3_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master onchip_memory2_3/s1 arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = onchip_memory2_3_s1_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master onchip_memory2_3/s1 arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = onchip_memory2_3_s1_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted onchip_memory2_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_3_s1 <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_3_s1 <= cpu_0_instruction_master_saved_grant_onchip_memory2_3_s1 ? 1 : (onchip_memory2_3_s1_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_onchip_memory2_3_s1) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_3_s1;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_0_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_0_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_0_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_0_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_0_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_0_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_0_instruction_master_requests_onchip_memory2_3_s1);

  //onchip_memory2_3_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign onchip_memory2_3_s1_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_0_instruction_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest;

  //cpu_1/data_master onchip_memory2_3/s1 arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = onchip_memory2_3_s1_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master onchip_memory2_3/s1 arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = onchip_memory2_3_s1_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted onchip_memory2_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_3_s1 <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_3_s1 <= cpu_1_data_master_saved_grant_onchip_memory2_3_s1 ? 1 : (onchip_memory2_3_s1_arbitration_holdoff_internal | ~cpu_1_data_master_requests_onchip_memory2_3_s1) ? 0 : last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_3_s1;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_3_s1 & cpu_1_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_3_s1 & cpu_1_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_3_s1 & cpu_1_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_3_s1 & cpu_1_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_3_s1 & cpu_1_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_3_s1 & cpu_1_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_data_master_granted_slave_onchip_memory2_3_s1 & cpu_1_data_master_requests_onchip_memory2_3_s1);

  //cpu_1/instruction_master onchip_memory2_3/s1 arbiterlock, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock = onchip_memory2_3_s1_slavearbiterlockenable & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master onchip_memory2_3/s1 arbiterlock2, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock2 = onchip_memory2_3_s1_slavearbiterlockenable2 & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master granted onchip_memory2_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_3_s1 <= 0;
      else 
        last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_3_s1 <= cpu_1_instruction_master_saved_grant_onchip_memory2_3_s1 ? 1 : (onchip_memory2_3_s1_arbitration_holdoff_internal | ~cpu_1_instruction_master_requests_onchip_memory2_3_s1) ? 0 : last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_3_s1;
    end


  //cpu_1_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_1_instruction_master_continuerequest = (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_1_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_1_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_1_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_1_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_1_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_1_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_1_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_1_instruction_master_requests_onchip_memory2_3_s1);

  //cpu_2/data_master onchip_memory2_3/s1 arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = onchip_memory2_3_s1_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master onchip_memory2_3/s1 arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = onchip_memory2_3_s1_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted onchip_memory2_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_3_s1 <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_3_s1 <= cpu_2_data_master_saved_grant_onchip_memory2_3_s1 ? 1 : (onchip_memory2_3_s1_arbitration_holdoff_internal | ~cpu_2_data_master_requests_onchip_memory2_3_s1) ? 0 : last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_3_s1;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_3_s1 & cpu_2_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_3_s1 & cpu_2_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_3_s1 & cpu_2_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_3_s1 & cpu_2_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_3_s1 & cpu_2_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_3_s1 & cpu_2_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_data_master_granted_slave_onchip_memory2_3_s1 & cpu_2_data_master_requests_onchip_memory2_3_s1);

  //cpu_2/instruction_master onchip_memory2_3/s1 arbiterlock, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock = onchip_memory2_3_s1_slavearbiterlockenable & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master onchip_memory2_3/s1 arbiterlock2, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock2 = onchip_memory2_3_s1_slavearbiterlockenable2 & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master granted onchip_memory2_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_3_s1 <= 0;
      else 
        last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_3_s1 <= cpu_2_instruction_master_saved_grant_onchip_memory2_3_s1 ? 1 : (onchip_memory2_3_s1_arbitration_holdoff_internal | ~cpu_2_instruction_master_requests_onchip_memory2_3_s1) ? 0 : last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_3_s1;
    end


  //cpu_2_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_2_instruction_master_continuerequest = (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_2_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_2_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_2_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_2_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_2_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_2_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_2_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_2_instruction_master_requests_onchip_memory2_3_s1);

  //cpu_3/data_master onchip_memory2_3/s1 arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = onchip_memory2_3_s1_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master onchip_memory2_3/s1 arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = onchip_memory2_3_s1_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted onchip_memory2_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_3_s1 <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_3_s1 <= cpu_3_data_master_saved_grant_onchip_memory2_3_s1 ? 1 : (onchip_memory2_3_s1_arbitration_holdoff_internal | ~cpu_3_data_master_requests_onchip_memory2_3_s1) ? 0 : last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_3_s1;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_3_s1 & cpu_3_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_3_s1 & cpu_3_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_3_s1 & cpu_3_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_3_s1 & cpu_3_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_3_s1 & cpu_3_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_3_s1 & cpu_3_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_data_master_granted_slave_onchip_memory2_3_s1 & cpu_3_data_master_requests_onchip_memory2_3_s1);

  //cpu_3/instruction_master onchip_memory2_3/s1 arbiterlock, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock = onchip_memory2_3_s1_slavearbiterlockenable & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master onchip_memory2_3/s1 arbiterlock2, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock2 = onchip_memory2_3_s1_slavearbiterlockenable2 & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master granted onchip_memory2_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_3_s1 <= 0;
      else 
        last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_3_s1 <= cpu_3_instruction_master_saved_grant_onchip_memory2_3_s1 ? 1 : (onchip_memory2_3_s1_arbitration_holdoff_internal | ~cpu_3_instruction_master_requests_onchip_memory2_3_s1) ? 0 : last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_3_s1;
    end


  //cpu_3_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_3_instruction_master_continuerequest = (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_3_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_3_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_3_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_3_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_3_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_3_instruction_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_3_instruction_master_granted_slave_onchip_memory2_3_s1 & cpu_3_instruction_master_requests_onchip_memory2_3_s1);

  assign cpu_0_data_master_qualified_request_onchip_memory2_3_s1 = cpu_0_data_master_requests_onchip_memory2_3_s1 & ~((cpu_0_data_master_read & ((1 < cpu_0_data_master_latency_counter) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in = cpu_0_data_master_granted_onchip_memory2_3_s1 & cpu_0_data_master_read & ~onchip_memory2_3_s1_waits_for_read;

  //shift register p1 cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register = {cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register, cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in};

  //cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register <= 0;
      else 
        cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register <= p1_cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
    end


  //local readdatavalid cpu_0_data_master_read_data_valid_onchip_memory2_3_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_onchip_memory2_3_s1 = cpu_0_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;

  //onchip_memory2_3_s1_writedata mux, which is an e_mux
  assign onchip_memory2_3_s1_writedata = (cpu_0_data_master_granted_onchip_memory2_3_s1)? cpu_0_data_master_writedata :
    (cpu_1_data_master_granted_onchip_memory2_3_s1)? cpu_1_data_master_writedata :
    (cpu_2_data_master_granted_onchip_memory2_3_s1)? cpu_2_data_master_writedata :
    cpu_3_data_master_writedata;

  //mux onchip_memory2_3_s1_clken, which is an e_mux
  assign onchip_memory2_3_s1_clken = 1'b1;

  assign cpu_0_instruction_master_requests_onchip_memory2_3_s1 = (({cpu_0_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h7000) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted onchip_memory2_3/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_3_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_3_s1 <= cpu_0_data_master_saved_grant_onchip_memory2_3_s1 ? 1 : (onchip_memory2_3_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_onchip_memory2_3_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_3_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_3_s1 & cpu_0_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_3_s1 & cpu_0_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_3_s1 & cpu_0_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_3_s1 & cpu_0_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_3_s1 & cpu_0_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_3_s1 & cpu_0_data_master_requests_onchip_memory2_3_s1) |
    (last_cycle_cpu_0_data_master_granted_slave_onchip_memory2_3_s1 & cpu_0_data_master_requests_onchip_memory2_3_s1);

  assign cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1 = cpu_0_instruction_master_requests_onchip_memory2_3_s1 & ~((cpu_0_instruction_master_read & ((1 < cpu_0_instruction_master_latency_counter))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in = cpu_0_instruction_master_granted_onchip_memory2_3_s1 & cpu_0_instruction_master_read & ~onchip_memory2_3_s1_waits_for_read;

  //shift register p1 cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register = {cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register, cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in};

  //cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register <= 0;
      else 
        cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register <= p1_cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
    end


  //local readdatavalid cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1 = cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;

  assign cpu_1_data_master_requests_onchip_memory2_3_s1 = ({cpu_1_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h7000) & (cpu_1_data_master_read | cpu_1_data_master_write);
  assign cpu_1_data_master_qualified_request_onchip_memory2_3_s1 = cpu_1_data_master_requests_onchip_memory2_3_s1 & ~((cpu_1_data_master_read & ((1 < cpu_1_data_master_latency_counter) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in = cpu_1_data_master_granted_onchip_memory2_3_s1 & cpu_1_data_master_read & ~onchip_memory2_3_s1_waits_for_read;

  //shift register p1 cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register = {cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register, cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in};

  //cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register <= 0;
      else 
        cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register <= p1_cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
    end


  //local readdatavalid cpu_1_data_master_read_data_valid_onchip_memory2_3_s1, which is an e_mux
  assign cpu_1_data_master_read_data_valid_onchip_memory2_3_s1 = cpu_1_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;

  assign cpu_1_instruction_master_requests_onchip_memory2_3_s1 = (({cpu_1_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h7000) & (cpu_1_instruction_master_read)) & cpu_1_instruction_master_read;
  assign cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1 = cpu_1_instruction_master_requests_onchip_memory2_3_s1 & ~((cpu_1_instruction_master_read & ((1 < cpu_1_instruction_master_latency_counter) | (|cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in = cpu_1_instruction_master_granted_onchip_memory2_3_s1 & cpu_1_instruction_master_read & ~onchip_memory2_3_s1_waits_for_read;

  //shift register p1 cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register = {cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register, cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in};

  //cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register <= 0;
      else 
        cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register <= p1_cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
    end


  //local readdatavalid cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1, which is an e_mux
  assign cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1 = cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;

  assign cpu_2_data_master_requests_onchip_memory2_3_s1 = ({cpu_2_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h7000) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_onchip_memory2_3_s1 = cpu_2_data_master_requests_onchip_memory2_3_s1 & ~((cpu_2_data_master_read & ((1 < cpu_2_data_master_latency_counter) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in = cpu_2_data_master_granted_onchip_memory2_3_s1 & cpu_2_data_master_read & ~onchip_memory2_3_s1_waits_for_read;

  //shift register p1 cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register = {cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register, cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in};

  //cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register <= 0;
      else 
        cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register <= p1_cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
    end


  //local readdatavalid cpu_2_data_master_read_data_valid_onchip_memory2_3_s1, which is an e_mux
  assign cpu_2_data_master_read_data_valid_onchip_memory2_3_s1 = cpu_2_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;

  assign cpu_2_instruction_master_requests_onchip_memory2_3_s1 = (({cpu_2_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h7000) & (cpu_2_instruction_master_read)) & cpu_2_instruction_master_read;
  assign cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1 = cpu_2_instruction_master_requests_onchip_memory2_3_s1 & ~((cpu_2_instruction_master_read & ((1 < cpu_2_instruction_master_latency_counter) | (|cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in = cpu_2_instruction_master_granted_onchip_memory2_3_s1 & cpu_2_instruction_master_read & ~onchip_memory2_3_s1_waits_for_read;

  //shift register p1 cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register = {cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register, cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in};

  //cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register <= 0;
      else 
        cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register <= p1_cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
    end


  //local readdatavalid cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1, which is an e_mux
  assign cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1 = cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;

  assign cpu_3_data_master_requests_onchip_memory2_3_s1 = ({cpu_3_data_master_address_to_slave[24 : 9] , 9'b0} == 25'h7000) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_onchip_memory2_3_s1 = cpu_3_data_master_requests_onchip_memory2_3_s1 & ~((cpu_3_data_master_read & ((1 < cpu_3_data_master_latency_counter) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in = cpu_3_data_master_granted_onchip_memory2_3_s1 & cpu_3_data_master_read & ~onchip_memory2_3_s1_waits_for_read;

  //shift register p1 cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register = {cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register, cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register_in};

  //cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register <= 0;
      else 
        cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register <= p1_cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;
    end


  //local readdatavalid cpu_3_data_master_read_data_valid_onchip_memory2_3_s1, which is an e_mux
  assign cpu_3_data_master_read_data_valid_onchip_memory2_3_s1 = cpu_3_data_master_read_data_valid_onchip_memory2_3_s1_shift_register;

  assign cpu_3_instruction_master_requests_onchip_memory2_3_s1 = (({cpu_3_instruction_master_address_to_slave[24 : 9] , 9'b0} == 25'h7000) & (cpu_3_instruction_master_read)) & cpu_3_instruction_master_read;
  assign cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1 = cpu_3_instruction_master_requests_onchip_memory2_3_s1 & ~((cpu_3_instruction_master_read & ((1 < cpu_3_instruction_master_latency_counter) | (|cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_0_instruction_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in = cpu_3_instruction_master_granted_onchip_memory2_3_s1 & cpu_3_instruction_master_read & ~onchip_memory2_3_s1_waits_for_read;

  //shift register p1 cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register = {cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register, cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register_in};

  //cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register <= 0;
      else 
        cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register <= p1_cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;
    end


  //local readdatavalid cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1, which is an e_mux
  assign cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1 = cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1_shift_register;

  //allow new arb cycle for onchip_memory2_3/s1, which is an e_assign
  assign onchip_memory2_3_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_1_instruction_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_2_instruction_master_arbiterlock & ~cpu_3_data_master_arbiterlock & ~cpu_3_instruction_master_arbiterlock;

  //cpu_3/instruction_master assignment into master qualified-requests vector for onchip_memory2_3/s1, which is an e_assign
  assign onchip_memory2_3_s1_master_qreq_vector[0] = cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1;

  //cpu_3/instruction_master grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_3_instruction_master_granted_onchip_memory2_3_s1 = onchip_memory2_3_s1_grant_vector[0];

  //cpu_3/instruction_master saved-grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_3_instruction_master_saved_grant_onchip_memory2_3_s1 = onchip_memory2_3_s1_arb_winner[0] && cpu_3_instruction_master_requests_onchip_memory2_3_s1;

  //cpu_3/data_master assignment into master qualified-requests vector for onchip_memory2_3/s1, which is an e_assign
  assign onchip_memory2_3_s1_master_qreq_vector[1] = cpu_3_data_master_qualified_request_onchip_memory2_3_s1;

  //cpu_3/data_master grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_3_data_master_granted_onchip_memory2_3_s1 = onchip_memory2_3_s1_grant_vector[1];

  //cpu_3/data_master saved-grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_3_data_master_saved_grant_onchip_memory2_3_s1 = onchip_memory2_3_s1_arb_winner[1] && cpu_3_data_master_requests_onchip_memory2_3_s1;

  //cpu_2/instruction_master assignment into master qualified-requests vector for onchip_memory2_3/s1, which is an e_assign
  assign onchip_memory2_3_s1_master_qreq_vector[2] = cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1;

  //cpu_2/instruction_master grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_2_instruction_master_granted_onchip_memory2_3_s1 = onchip_memory2_3_s1_grant_vector[2];

  //cpu_2/instruction_master saved-grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_2_instruction_master_saved_grant_onchip_memory2_3_s1 = onchip_memory2_3_s1_arb_winner[2] && cpu_2_instruction_master_requests_onchip_memory2_3_s1;

  //cpu_2/data_master assignment into master qualified-requests vector for onchip_memory2_3/s1, which is an e_assign
  assign onchip_memory2_3_s1_master_qreq_vector[3] = cpu_2_data_master_qualified_request_onchip_memory2_3_s1;

  //cpu_2/data_master grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_2_data_master_granted_onchip_memory2_3_s1 = onchip_memory2_3_s1_grant_vector[3];

  //cpu_2/data_master saved-grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_2_data_master_saved_grant_onchip_memory2_3_s1 = onchip_memory2_3_s1_arb_winner[3] && cpu_2_data_master_requests_onchip_memory2_3_s1;

  //cpu_1/instruction_master assignment into master qualified-requests vector for onchip_memory2_3/s1, which is an e_assign
  assign onchip_memory2_3_s1_master_qreq_vector[4] = cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1;

  //cpu_1/instruction_master grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_1_instruction_master_granted_onchip_memory2_3_s1 = onchip_memory2_3_s1_grant_vector[4];

  //cpu_1/instruction_master saved-grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_1_instruction_master_saved_grant_onchip_memory2_3_s1 = onchip_memory2_3_s1_arb_winner[4] && cpu_1_instruction_master_requests_onchip_memory2_3_s1;

  //cpu_1/data_master assignment into master qualified-requests vector for onchip_memory2_3/s1, which is an e_assign
  assign onchip_memory2_3_s1_master_qreq_vector[5] = cpu_1_data_master_qualified_request_onchip_memory2_3_s1;

  //cpu_1/data_master grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_1_data_master_granted_onchip_memory2_3_s1 = onchip_memory2_3_s1_grant_vector[5];

  //cpu_1/data_master saved-grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_1_data_master_saved_grant_onchip_memory2_3_s1 = onchip_memory2_3_s1_arb_winner[5] && cpu_1_data_master_requests_onchip_memory2_3_s1;

  //cpu_0/instruction_master assignment into master qualified-requests vector for onchip_memory2_3/s1, which is an e_assign
  assign onchip_memory2_3_s1_master_qreq_vector[6] = cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1;

  //cpu_0/instruction_master grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_0_instruction_master_granted_onchip_memory2_3_s1 = onchip_memory2_3_s1_grant_vector[6];

  //cpu_0/instruction_master saved-grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_onchip_memory2_3_s1 = onchip_memory2_3_s1_arb_winner[6] && cpu_0_instruction_master_requests_onchip_memory2_3_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for onchip_memory2_3/s1, which is an e_assign
  assign onchip_memory2_3_s1_master_qreq_vector[7] = cpu_0_data_master_qualified_request_onchip_memory2_3_s1;

  //cpu_0/data_master grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_0_data_master_granted_onchip_memory2_3_s1 = onchip_memory2_3_s1_grant_vector[7];

  //cpu_0/data_master saved-grant onchip_memory2_3/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_onchip_memory2_3_s1 = onchip_memory2_3_s1_arb_winner[7] && cpu_0_data_master_requests_onchip_memory2_3_s1;

  //onchip_memory2_3/s1 chosen-master double-vector, which is an e_assign
  assign onchip_memory2_3_s1_chosen_master_double_vector = {onchip_memory2_3_s1_master_qreq_vector, onchip_memory2_3_s1_master_qreq_vector} & ({~onchip_memory2_3_s1_master_qreq_vector, ~onchip_memory2_3_s1_master_qreq_vector} + onchip_memory2_3_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign onchip_memory2_3_s1_arb_winner = (onchip_memory2_3_s1_allow_new_arb_cycle & | onchip_memory2_3_s1_grant_vector) ? onchip_memory2_3_s1_grant_vector : onchip_memory2_3_s1_saved_chosen_master_vector;

  //saved onchip_memory2_3_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_3_s1_saved_chosen_master_vector <= 0;
      else if (onchip_memory2_3_s1_allow_new_arb_cycle)
          onchip_memory2_3_s1_saved_chosen_master_vector <= |onchip_memory2_3_s1_grant_vector ? onchip_memory2_3_s1_grant_vector : onchip_memory2_3_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign onchip_memory2_3_s1_grant_vector = {(onchip_memory2_3_s1_chosen_master_double_vector[7] | onchip_memory2_3_s1_chosen_master_double_vector[15]),
    (onchip_memory2_3_s1_chosen_master_double_vector[6] | onchip_memory2_3_s1_chosen_master_double_vector[14]),
    (onchip_memory2_3_s1_chosen_master_double_vector[5] | onchip_memory2_3_s1_chosen_master_double_vector[13]),
    (onchip_memory2_3_s1_chosen_master_double_vector[4] | onchip_memory2_3_s1_chosen_master_double_vector[12]),
    (onchip_memory2_3_s1_chosen_master_double_vector[3] | onchip_memory2_3_s1_chosen_master_double_vector[11]),
    (onchip_memory2_3_s1_chosen_master_double_vector[2] | onchip_memory2_3_s1_chosen_master_double_vector[10]),
    (onchip_memory2_3_s1_chosen_master_double_vector[1] | onchip_memory2_3_s1_chosen_master_double_vector[9]),
    (onchip_memory2_3_s1_chosen_master_double_vector[0] | onchip_memory2_3_s1_chosen_master_double_vector[8])};

  //onchip_memory2_3/s1 chosen master rotated left, which is an e_assign
  assign onchip_memory2_3_s1_chosen_master_rot_left = (onchip_memory2_3_s1_arb_winner << 1) ? (onchip_memory2_3_s1_arb_winner << 1) : 1;

  //onchip_memory2_3/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_3_s1_arb_addend <= 1;
      else if (|onchip_memory2_3_s1_grant_vector)
          onchip_memory2_3_s1_arb_addend <= onchip_memory2_3_s1_end_xfer? onchip_memory2_3_s1_chosen_master_rot_left : onchip_memory2_3_s1_grant_vector;
    end


  //~onchip_memory2_3_s1_reset assignment, which is an e_assign
  assign onchip_memory2_3_s1_reset = ~reset_n;

  assign onchip_memory2_3_s1_chipselect = cpu_0_data_master_granted_onchip_memory2_3_s1 | cpu_0_instruction_master_granted_onchip_memory2_3_s1 | cpu_1_data_master_granted_onchip_memory2_3_s1 | cpu_1_instruction_master_granted_onchip_memory2_3_s1 | cpu_2_data_master_granted_onchip_memory2_3_s1 | cpu_2_instruction_master_granted_onchip_memory2_3_s1 | cpu_3_data_master_granted_onchip_memory2_3_s1 | cpu_3_instruction_master_granted_onchip_memory2_3_s1;
  //onchip_memory2_3_s1_firsttransfer first transaction, which is an e_assign
  assign onchip_memory2_3_s1_firsttransfer = onchip_memory2_3_s1_begins_xfer ? onchip_memory2_3_s1_unreg_firsttransfer : onchip_memory2_3_s1_reg_firsttransfer;

  //onchip_memory2_3_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign onchip_memory2_3_s1_unreg_firsttransfer = ~(onchip_memory2_3_s1_slavearbiterlockenable & onchip_memory2_3_s1_any_continuerequest);

  //onchip_memory2_3_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          onchip_memory2_3_s1_reg_firsttransfer <= 1'b1;
      else if (onchip_memory2_3_s1_begins_xfer)
          onchip_memory2_3_s1_reg_firsttransfer <= onchip_memory2_3_s1_unreg_firsttransfer;
    end


  //onchip_memory2_3_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign onchip_memory2_3_s1_beginbursttransfer_internal = onchip_memory2_3_s1_begins_xfer;

  //onchip_memory2_3_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign onchip_memory2_3_s1_arbitration_holdoff_internal = onchip_memory2_3_s1_begins_xfer & onchip_memory2_3_s1_firsttransfer;

  //onchip_memory2_3_s1_write assignment, which is an e_mux
  assign onchip_memory2_3_s1_write = (cpu_0_data_master_granted_onchip_memory2_3_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_onchip_memory2_3_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_onchip_memory2_3_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_onchip_memory2_3_s1 & cpu_3_data_master_write);

  assign shifted_address_to_onchip_memory2_3_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //onchip_memory2_3_s1_address mux, which is an e_mux
  assign onchip_memory2_3_s1_address = (cpu_0_data_master_granted_onchip_memory2_3_s1)? (shifted_address_to_onchip_memory2_3_s1_from_cpu_0_data_master >> 2) :
    (cpu_0_instruction_master_granted_onchip_memory2_3_s1)? (shifted_address_to_onchip_memory2_3_s1_from_cpu_0_instruction_master >> 2) :
    (cpu_1_data_master_granted_onchip_memory2_3_s1)? (shifted_address_to_onchip_memory2_3_s1_from_cpu_1_data_master >> 2) :
    (cpu_1_instruction_master_granted_onchip_memory2_3_s1)? (shifted_address_to_onchip_memory2_3_s1_from_cpu_1_instruction_master >> 2) :
    (cpu_2_data_master_granted_onchip_memory2_3_s1)? (shifted_address_to_onchip_memory2_3_s1_from_cpu_2_data_master >> 2) :
    (cpu_2_instruction_master_granted_onchip_memory2_3_s1)? (shifted_address_to_onchip_memory2_3_s1_from_cpu_2_instruction_master >> 2) :
    (cpu_3_data_master_granted_onchip_memory2_3_s1)? (shifted_address_to_onchip_memory2_3_s1_from_cpu_3_data_master >> 2) :
    (shifted_address_to_onchip_memory2_3_s1_from_cpu_3_instruction_master >> 2);

  assign shifted_address_to_onchip_memory2_3_s1_from_cpu_0_instruction_master = cpu_0_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_3_s1_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_3_s1_from_cpu_1_instruction_master = cpu_1_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_3_s1_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_3_s1_from_cpu_2_instruction_master = cpu_2_instruction_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_3_s1_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  assign shifted_address_to_onchip_memory2_3_s1_from_cpu_3_instruction_master = cpu_3_instruction_master_address_to_slave;
  //d1_onchip_memory2_3_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_onchip_memory2_3_s1_end_xfer <= 1;
      else 
        d1_onchip_memory2_3_s1_end_xfer <= onchip_memory2_3_s1_end_xfer;
    end


  //onchip_memory2_3_s1_waits_for_read in a cycle, which is an e_mux
  assign onchip_memory2_3_s1_waits_for_read = onchip_memory2_3_s1_in_a_read_cycle & 0;

  //onchip_memory2_3_s1_in_a_read_cycle assignment, which is an e_assign
  assign onchip_memory2_3_s1_in_a_read_cycle = (cpu_0_data_master_granted_onchip_memory2_3_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_onchip_memory2_3_s1 & cpu_0_instruction_master_read) | (cpu_1_data_master_granted_onchip_memory2_3_s1 & cpu_1_data_master_read) | (cpu_1_instruction_master_granted_onchip_memory2_3_s1 & cpu_1_instruction_master_read) | (cpu_2_data_master_granted_onchip_memory2_3_s1 & cpu_2_data_master_read) | (cpu_2_instruction_master_granted_onchip_memory2_3_s1 & cpu_2_instruction_master_read) | (cpu_3_data_master_granted_onchip_memory2_3_s1 & cpu_3_data_master_read) | (cpu_3_instruction_master_granted_onchip_memory2_3_s1 & cpu_3_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = onchip_memory2_3_s1_in_a_read_cycle;

  //onchip_memory2_3_s1_waits_for_write in a cycle, which is an e_mux
  assign onchip_memory2_3_s1_waits_for_write = onchip_memory2_3_s1_in_a_write_cycle & 0;

  //onchip_memory2_3_s1_in_a_write_cycle assignment, which is an e_assign
  assign onchip_memory2_3_s1_in_a_write_cycle = (cpu_0_data_master_granted_onchip_memory2_3_s1 & cpu_0_data_master_write) | (cpu_1_data_master_granted_onchip_memory2_3_s1 & cpu_1_data_master_write) | (cpu_2_data_master_granted_onchip_memory2_3_s1 & cpu_2_data_master_write) | (cpu_3_data_master_granted_onchip_memory2_3_s1 & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = onchip_memory2_3_s1_in_a_write_cycle;

  assign wait_for_onchip_memory2_3_s1_counter = 0;
  //onchip_memory2_3_s1_byteenable byte enable port mux, which is an e_mux
  assign onchip_memory2_3_s1_byteenable = (cpu_0_data_master_granted_onchip_memory2_3_s1)? cpu_0_data_master_byteenable :
    (cpu_1_data_master_granted_onchip_memory2_3_s1)? cpu_1_data_master_byteenable :
    (cpu_2_data_master_granted_onchip_memory2_3_s1)? cpu_2_data_master_byteenable :
    (cpu_3_data_master_granted_onchip_memory2_3_s1)? cpu_3_data_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //onchip_memory2_3/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_onchip_memory2_3_s1 + cpu_0_instruction_master_granted_onchip_memory2_3_s1 + cpu_1_data_master_granted_onchip_memory2_3_s1 + cpu_1_instruction_master_granted_onchip_memory2_3_s1 + cpu_2_data_master_granted_onchip_memory2_3_s1 + cpu_2_instruction_master_granted_onchip_memory2_3_s1 + cpu_3_data_master_granted_onchip_memory2_3_s1 + cpu_3_instruction_master_granted_onchip_memory2_3_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_onchip_memory2_3_s1 + cpu_0_instruction_master_saved_grant_onchip_memory2_3_s1 + cpu_1_data_master_saved_grant_onchip_memory2_3_s1 + cpu_1_instruction_master_saved_grant_onchip_memory2_3_s1 + cpu_2_data_master_saved_grant_onchip_memory2_3_s1 + cpu_2_instruction_master_saved_grant_onchip_memory2_3_s1 + cpu_3_data_master_saved_grant_onchip_memory2_3_s1 + cpu_3_instruction_master_saved_grant_onchip_memory2_3_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module performance_counter_0_control_slave_arbitrator (
                                                        // inputs:
                                                         clk,
                                                         cpu_0_data_master_address_to_slave,
                                                         cpu_0_data_master_latency_counter,
                                                         cpu_0_data_master_read,
                                                         cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                         cpu_0_data_master_write,
                                                         cpu_0_data_master_writedata,
                                                         cpu_1_data_master_address_to_slave,
                                                         cpu_1_data_master_latency_counter,
                                                         cpu_1_data_master_read,
                                                         cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                         cpu_1_data_master_write,
                                                         cpu_1_data_master_writedata,
                                                         cpu_2_data_master_address_to_slave,
                                                         cpu_2_data_master_latency_counter,
                                                         cpu_2_data_master_read,
                                                         cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                         cpu_2_data_master_write,
                                                         cpu_2_data_master_writedata,
                                                         cpu_3_data_master_address_to_slave,
                                                         cpu_3_data_master_latency_counter,
                                                         cpu_3_data_master_read,
                                                         cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                         cpu_3_data_master_write,
                                                         cpu_3_data_master_writedata,
                                                         performance_counter_0_control_slave_readdata,
                                                         reset_n,

                                                        // outputs:
                                                         cpu_0_data_master_granted_performance_counter_0_control_slave,
                                                         cpu_0_data_master_qualified_request_performance_counter_0_control_slave,
                                                         cpu_0_data_master_read_data_valid_performance_counter_0_control_slave,
                                                         cpu_0_data_master_requests_performance_counter_0_control_slave,
                                                         cpu_1_data_master_granted_performance_counter_0_control_slave,
                                                         cpu_1_data_master_qualified_request_performance_counter_0_control_slave,
                                                         cpu_1_data_master_read_data_valid_performance_counter_0_control_slave,
                                                         cpu_1_data_master_requests_performance_counter_0_control_slave,
                                                         cpu_2_data_master_granted_performance_counter_0_control_slave,
                                                         cpu_2_data_master_qualified_request_performance_counter_0_control_slave,
                                                         cpu_2_data_master_read_data_valid_performance_counter_0_control_slave,
                                                         cpu_2_data_master_requests_performance_counter_0_control_slave,
                                                         cpu_3_data_master_granted_performance_counter_0_control_slave,
                                                         cpu_3_data_master_qualified_request_performance_counter_0_control_slave,
                                                         cpu_3_data_master_read_data_valid_performance_counter_0_control_slave,
                                                         cpu_3_data_master_requests_performance_counter_0_control_slave,
                                                         d1_performance_counter_0_control_slave_end_xfer,
                                                         performance_counter_0_control_slave_address,
                                                         performance_counter_0_control_slave_begintransfer,
                                                         performance_counter_0_control_slave_readdata_from_sa,
                                                         performance_counter_0_control_slave_reset_n,
                                                         performance_counter_0_control_slave_write,
                                                         performance_counter_0_control_slave_writedata
                                                      )
;

  output           cpu_0_data_master_granted_performance_counter_0_control_slave;
  output           cpu_0_data_master_qualified_request_performance_counter_0_control_slave;
  output           cpu_0_data_master_read_data_valid_performance_counter_0_control_slave;
  output           cpu_0_data_master_requests_performance_counter_0_control_slave;
  output           cpu_1_data_master_granted_performance_counter_0_control_slave;
  output           cpu_1_data_master_qualified_request_performance_counter_0_control_slave;
  output           cpu_1_data_master_read_data_valid_performance_counter_0_control_slave;
  output           cpu_1_data_master_requests_performance_counter_0_control_slave;
  output           cpu_2_data_master_granted_performance_counter_0_control_slave;
  output           cpu_2_data_master_qualified_request_performance_counter_0_control_slave;
  output           cpu_2_data_master_read_data_valid_performance_counter_0_control_slave;
  output           cpu_2_data_master_requests_performance_counter_0_control_slave;
  output           cpu_3_data_master_granted_performance_counter_0_control_slave;
  output           cpu_3_data_master_qualified_request_performance_counter_0_control_slave;
  output           cpu_3_data_master_read_data_valid_performance_counter_0_control_slave;
  output           cpu_3_data_master_requests_performance_counter_0_control_slave;
  output           d1_performance_counter_0_control_slave_end_xfer;
  output  [  3: 0] performance_counter_0_control_slave_address;
  output           performance_counter_0_control_slave_begintransfer;
  output  [ 31: 0] performance_counter_0_control_slave_readdata_from_sa;
  output           performance_counter_0_control_slave_reset_n;
  output           performance_counter_0_control_slave_write;
  output  [ 31: 0] performance_counter_0_control_slave_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input   [ 31: 0] performance_counter_0_control_slave_readdata;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_performance_counter_0_control_slave;
  wire             cpu_0_data_master_qualified_request_performance_counter_0_control_slave;
  wire             cpu_0_data_master_read_data_valid_performance_counter_0_control_slave;
  reg              cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
  wire             cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in;
  wire             cpu_0_data_master_requests_performance_counter_0_control_slave;
  wire             cpu_0_data_master_saved_grant_performance_counter_0_control_slave;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_performance_counter_0_control_slave;
  wire             cpu_1_data_master_qualified_request_performance_counter_0_control_slave;
  wire             cpu_1_data_master_read_data_valid_performance_counter_0_control_slave;
  reg              cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
  wire             cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in;
  wire             cpu_1_data_master_requests_performance_counter_0_control_slave;
  wire             cpu_1_data_master_saved_grant_performance_counter_0_control_slave;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_performance_counter_0_control_slave;
  wire             cpu_2_data_master_qualified_request_performance_counter_0_control_slave;
  wire             cpu_2_data_master_read_data_valid_performance_counter_0_control_slave;
  reg              cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
  wire             cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in;
  wire             cpu_2_data_master_requests_performance_counter_0_control_slave;
  wire             cpu_2_data_master_saved_grant_performance_counter_0_control_slave;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_performance_counter_0_control_slave;
  wire             cpu_3_data_master_qualified_request_performance_counter_0_control_slave;
  wire             cpu_3_data_master_read_data_valid_performance_counter_0_control_slave;
  reg              cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
  wire             cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in;
  wire             cpu_3_data_master_requests_performance_counter_0_control_slave;
  wire             cpu_3_data_master_saved_grant_performance_counter_0_control_slave;
  reg              d1_performance_counter_0_control_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_performance_counter_0_control_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_performance_counter_0_control_slave;
  reg              last_cycle_cpu_1_data_master_granted_slave_performance_counter_0_control_slave;
  reg              last_cycle_cpu_2_data_master_granted_slave_performance_counter_0_control_slave;
  reg              last_cycle_cpu_3_data_master_granted_slave_performance_counter_0_control_slave;
  wire             p1_cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
  wire             p1_cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
  wire             p1_cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
  wire             p1_cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
  wire    [  3: 0] performance_counter_0_control_slave_address;
  wire             performance_counter_0_control_slave_allgrants;
  wire             performance_counter_0_control_slave_allow_new_arb_cycle;
  wire             performance_counter_0_control_slave_any_bursting_master_saved_grant;
  wire             performance_counter_0_control_slave_any_continuerequest;
  reg     [  3: 0] performance_counter_0_control_slave_arb_addend;
  wire             performance_counter_0_control_slave_arb_counter_enable;
  reg     [  2: 0] performance_counter_0_control_slave_arb_share_counter;
  wire    [  2: 0] performance_counter_0_control_slave_arb_share_counter_next_value;
  wire    [  2: 0] performance_counter_0_control_slave_arb_share_set_values;
  wire    [  3: 0] performance_counter_0_control_slave_arb_winner;
  wire             performance_counter_0_control_slave_arbitration_holdoff_internal;
  wire             performance_counter_0_control_slave_beginbursttransfer_internal;
  wire             performance_counter_0_control_slave_begins_xfer;
  wire             performance_counter_0_control_slave_begintransfer;
  wire    [  7: 0] performance_counter_0_control_slave_chosen_master_double_vector;
  wire    [  3: 0] performance_counter_0_control_slave_chosen_master_rot_left;
  wire             performance_counter_0_control_slave_end_xfer;
  wire             performance_counter_0_control_slave_firsttransfer;
  wire    [  3: 0] performance_counter_0_control_slave_grant_vector;
  wire             performance_counter_0_control_slave_in_a_read_cycle;
  wire             performance_counter_0_control_slave_in_a_write_cycle;
  wire    [  3: 0] performance_counter_0_control_slave_master_qreq_vector;
  wire             performance_counter_0_control_slave_non_bursting_master_requests;
  wire    [ 31: 0] performance_counter_0_control_slave_readdata_from_sa;
  reg              performance_counter_0_control_slave_reg_firsttransfer;
  wire             performance_counter_0_control_slave_reset_n;
  reg     [  3: 0] performance_counter_0_control_slave_saved_chosen_master_vector;
  reg              performance_counter_0_control_slave_slavearbiterlockenable;
  wire             performance_counter_0_control_slave_slavearbiterlockenable2;
  wire             performance_counter_0_control_slave_unreg_firsttransfer;
  wire             performance_counter_0_control_slave_waits_for_read;
  wire             performance_counter_0_control_slave_waits_for_write;
  wire             performance_counter_0_control_slave_write;
  wire    [ 31: 0] performance_counter_0_control_slave_writedata;
  wire    [ 24: 0] shifted_address_to_performance_counter_0_control_slave_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_performance_counter_0_control_slave_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_performance_counter_0_control_slave_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_performance_counter_0_control_slave_from_cpu_3_data_master;
  wire             wait_for_performance_counter_0_control_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~performance_counter_0_control_slave_end_xfer;
    end


  assign performance_counter_0_control_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_performance_counter_0_control_slave | cpu_1_data_master_qualified_request_performance_counter_0_control_slave | cpu_2_data_master_qualified_request_performance_counter_0_control_slave | cpu_3_data_master_qualified_request_performance_counter_0_control_slave));
  //assign performance_counter_0_control_slave_readdata_from_sa = performance_counter_0_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign performance_counter_0_control_slave_readdata_from_sa = performance_counter_0_control_slave_readdata;

  assign cpu_0_data_master_requests_performance_counter_0_control_slave = ({cpu_0_data_master_address_to_slave[24 : 6] , 6'b0} == 25'h0) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //performance_counter_0_control_slave_arb_share_counter set values, which is an e_mux
  assign performance_counter_0_control_slave_arb_share_set_values = 1;

  //performance_counter_0_control_slave_non_bursting_master_requests mux, which is an e_mux
  assign performance_counter_0_control_slave_non_bursting_master_requests = cpu_0_data_master_requests_performance_counter_0_control_slave |
    cpu_1_data_master_requests_performance_counter_0_control_slave |
    cpu_2_data_master_requests_performance_counter_0_control_slave |
    cpu_3_data_master_requests_performance_counter_0_control_slave |
    cpu_0_data_master_requests_performance_counter_0_control_slave |
    cpu_1_data_master_requests_performance_counter_0_control_slave |
    cpu_2_data_master_requests_performance_counter_0_control_slave |
    cpu_3_data_master_requests_performance_counter_0_control_slave |
    cpu_0_data_master_requests_performance_counter_0_control_slave |
    cpu_1_data_master_requests_performance_counter_0_control_slave |
    cpu_2_data_master_requests_performance_counter_0_control_slave |
    cpu_3_data_master_requests_performance_counter_0_control_slave |
    cpu_0_data_master_requests_performance_counter_0_control_slave |
    cpu_1_data_master_requests_performance_counter_0_control_slave |
    cpu_2_data_master_requests_performance_counter_0_control_slave |
    cpu_3_data_master_requests_performance_counter_0_control_slave;

  //performance_counter_0_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign performance_counter_0_control_slave_any_bursting_master_saved_grant = 0;

  //performance_counter_0_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign performance_counter_0_control_slave_arb_share_counter_next_value = performance_counter_0_control_slave_firsttransfer ? (performance_counter_0_control_slave_arb_share_set_values - 1) : |performance_counter_0_control_slave_arb_share_counter ? (performance_counter_0_control_slave_arb_share_counter - 1) : 0;

  //performance_counter_0_control_slave_allgrants all slave grants, which is an e_mux
  assign performance_counter_0_control_slave_allgrants = (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector) |
    (|performance_counter_0_control_slave_grant_vector);

  //performance_counter_0_control_slave_end_xfer assignment, which is an e_assign
  assign performance_counter_0_control_slave_end_xfer = ~(performance_counter_0_control_slave_waits_for_read | performance_counter_0_control_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_performance_counter_0_control_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_performance_counter_0_control_slave = performance_counter_0_control_slave_end_xfer & (~performance_counter_0_control_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //performance_counter_0_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign performance_counter_0_control_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_performance_counter_0_control_slave & performance_counter_0_control_slave_allgrants) | (end_xfer_arb_share_counter_term_performance_counter_0_control_slave & ~performance_counter_0_control_slave_non_bursting_master_requests);

  //performance_counter_0_control_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          performance_counter_0_control_slave_arb_share_counter <= 0;
      else if (performance_counter_0_control_slave_arb_counter_enable)
          performance_counter_0_control_slave_arb_share_counter <= performance_counter_0_control_slave_arb_share_counter_next_value;
    end


  //performance_counter_0_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          performance_counter_0_control_slave_slavearbiterlockenable <= 0;
      else if ((|performance_counter_0_control_slave_master_qreq_vector & end_xfer_arb_share_counter_term_performance_counter_0_control_slave) | (end_xfer_arb_share_counter_term_performance_counter_0_control_slave & ~performance_counter_0_control_slave_non_bursting_master_requests))
          performance_counter_0_control_slave_slavearbiterlockenable <= |performance_counter_0_control_slave_arb_share_counter_next_value;
    end


  //cpu_0/data_master performance_counter_0/control_slave arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = performance_counter_0_control_slave_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //performance_counter_0_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign performance_counter_0_control_slave_slavearbiterlockenable2 = |performance_counter_0_control_slave_arb_share_counter_next_value;

  //cpu_0/data_master performance_counter_0/control_slave arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = performance_counter_0_control_slave_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_1/data_master performance_counter_0/control_slave arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = performance_counter_0_control_slave_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master performance_counter_0/control_slave arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = performance_counter_0_control_slave_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted performance_counter_0/control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_performance_counter_0_control_slave <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_performance_counter_0_control_slave <= cpu_1_data_master_saved_grant_performance_counter_0_control_slave ? 1 : (performance_counter_0_control_slave_arbitration_holdoff_internal | ~cpu_1_data_master_requests_performance_counter_0_control_slave) ? 0 : last_cycle_cpu_1_data_master_granted_slave_performance_counter_0_control_slave;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_performance_counter_0_control_slave & cpu_1_data_master_requests_performance_counter_0_control_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_performance_counter_0_control_slave & cpu_1_data_master_requests_performance_counter_0_control_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_performance_counter_0_control_slave & cpu_1_data_master_requests_performance_counter_0_control_slave);

  //performance_counter_0_control_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  assign performance_counter_0_control_slave_any_continuerequest = cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest;

  //cpu_2/data_master performance_counter_0/control_slave arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = performance_counter_0_control_slave_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master performance_counter_0/control_slave arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = performance_counter_0_control_slave_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted performance_counter_0/control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_performance_counter_0_control_slave <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_performance_counter_0_control_slave <= cpu_2_data_master_saved_grant_performance_counter_0_control_slave ? 1 : (performance_counter_0_control_slave_arbitration_holdoff_internal | ~cpu_2_data_master_requests_performance_counter_0_control_slave) ? 0 : last_cycle_cpu_2_data_master_granted_slave_performance_counter_0_control_slave;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_performance_counter_0_control_slave & cpu_2_data_master_requests_performance_counter_0_control_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_performance_counter_0_control_slave & cpu_2_data_master_requests_performance_counter_0_control_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_performance_counter_0_control_slave & cpu_2_data_master_requests_performance_counter_0_control_slave);

  //cpu_3/data_master performance_counter_0/control_slave arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = performance_counter_0_control_slave_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master performance_counter_0/control_slave arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = performance_counter_0_control_slave_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted performance_counter_0/control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_performance_counter_0_control_slave <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_performance_counter_0_control_slave <= cpu_3_data_master_saved_grant_performance_counter_0_control_slave ? 1 : (performance_counter_0_control_slave_arbitration_holdoff_internal | ~cpu_3_data_master_requests_performance_counter_0_control_slave) ? 0 : last_cycle_cpu_3_data_master_granted_slave_performance_counter_0_control_slave;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_performance_counter_0_control_slave & cpu_3_data_master_requests_performance_counter_0_control_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_performance_counter_0_control_slave & cpu_3_data_master_requests_performance_counter_0_control_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_performance_counter_0_control_slave & cpu_3_data_master_requests_performance_counter_0_control_slave);

  assign cpu_0_data_master_qualified_request_performance_counter_0_control_slave = cpu_0_data_master_requests_performance_counter_0_control_slave & ~((cpu_0_data_master_read & ((1 < cpu_0_data_master_latency_counter) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in = cpu_0_data_master_granted_performance_counter_0_control_slave & cpu_0_data_master_read & ~performance_counter_0_control_slave_waits_for_read;

  //shift register p1 cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register = {cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register, cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in};

  //cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register <= 0;
      else 
        cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register <= p1_cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
    end


  //local readdatavalid cpu_0_data_master_read_data_valid_performance_counter_0_control_slave, which is an e_mux
  assign cpu_0_data_master_read_data_valid_performance_counter_0_control_slave = cpu_0_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;

  //performance_counter_0_control_slave_writedata mux, which is an e_mux
  assign performance_counter_0_control_slave_writedata = (cpu_0_data_master_granted_performance_counter_0_control_slave)? cpu_0_data_master_writedata :
    (cpu_1_data_master_granted_performance_counter_0_control_slave)? cpu_1_data_master_writedata :
    (cpu_2_data_master_granted_performance_counter_0_control_slave)? cpu_2_data_master_writedata :
    cpu_3_data_master_writedata;

  assign cpu_1_data_master_requests_performance_counter_0_control_slave = ({cpu_1_data_master_address_to_slave[24 : 6] , 6'b0} == 25'h0) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //cpu_0/data_master granted performance_counter_0/control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_performance_counter_0_control_slave <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_performance_counter_0_control_slave <= cpu_0_data_master_saved_grant_performance_counter_0_control_slave ? 1 : (performance_counter_0_control_slave_arbitration_holdoff_internal | ~cpu_0_data_master_requests_performance_counter_0_control_slave) ? 0 : last_cycle_cpu_0_data_master_granted_slave_performance_counter_0_control_slave;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_performance_counter_0_control_slave & cpu_0_data_master_requests_performance_counter_0_control_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_performance_counter_0_control_slave & cpu_0_data_master_requests_performance_counter_0_control_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_performance_counter_0_control_slave & cpu_0_data_master_requests_performance_counter_0_control_slave);

  assign cpu_1_data_master_qualified_request_performance_counter_0_control_slave = cpu_1_data_master_requests_performance_counter_0_control_slave & ~((cpu_1_data_master_read & ((1 < cpu_1_data_master_latency_counter) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in = cpu_1_data_master_granted_performance_counter_0_control_slave & cpu_1_data_master_read & ~performance_counter_0_control_slave_waits_for_read;

  //shift register p1 cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register = {cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register, cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in};

  //cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register <= 0;
      else 
        cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register <= p1_cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
    end


  //local readdatavalid cpu_1_data_master_read_data_valid_performance_counter_0_control_slave, which is an e_mux
  assign cpu_1_data_master_read_data_valid_performance_counter_0_control_slave = cpu_1_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;

  assign cpu_2_data_master_requests_performance_counter_0_control_slave = ({cpu_2_data_master_address_to_slave[24 : 6] , 6'b0} == 25'h0) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_performance_counter_0_control_slave = cpu_2_data_master_requests_performance_counter_0_control_slave & ~((cpu_2_data_master_read & ((1 < cpu_2_data_master_latency_counter) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in = cpu_2_data_master_granted_performance_counter_0_control_slave & cpu_2_data_master_read & ~performance_counter_0_control_slave_waits_for_read;

  //shift register p1 cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register = {cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register, cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in};

  //cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register <= 0;
      else 
        cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register <= p1_cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
    end


  //local readdatavalid cpu_2_data_master_read_data_valid_performance_counter_0_control_slave, which is an e_mux
  assign cpu_2_data_master_read_data_valid_performance_counter_0_control_slave = cpu_2_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;

  assign cpu_3_data_master_requests_performance_counter_0_control_slave = ({cpu_3_data_master_address_to_slave[24 : 6] , 6'b0} == 25'h0) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_performance_counter_0_control_slave = cpu_3_data_master_requests_performance_counter_0_control_slave & ~((cpu_3_data_master_read & ((1 < cpu_3_data_master_latency_counter) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock);
  //cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in = cpu_3_data_master_granted_performance_counter_0_control_slave & cpu_3_data_master_read & ~performance_counter_0_control_slave_waits_for_read;

  //shift register p1 cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register = {cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register, cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register_in};

  //cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register <= 0;
      else 
        cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register <= p1_cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;
    end


  //local readdatavalid cpu_3_data_master_read_data_valid_performance_counter_0_control_slave, which is an e_mux
  assign cpu_3_data_master_read_data_valid_performance_counter_0_control_slave = cpu_3_data_master_read_data_valid_performance_counter_0_control_slave_shift_register;

  //allow new arb cycle for performance_counter_0/control_slave, which is an e_assign
  assign performance_counter_0_control_slave_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_3_data_master_arbiterlock;

  //cpu_3/data_master assignment into master qualified-requests vector for performance_counter_0/control_slave, which is an e_assign
  assign performance_counter_0_control_slave_master_qreq_vector[0] = cpu_3_data_master_qualified_request_performance_counter_0_control_slave;

  //cpu_3/data_master grant performance_counter_0/control_slave, which is an e_assign
  assign cpu_3_data_master_granted_performance_counter_0_control_slave = performance_counter_0_control_slave_grant_vector[0];

  //cpu_3/data_master saved-grant performance_counter_0/control_slave, which is an e_assign
  assign cpu_3_data_master_saved_grant_performance_counter_0_control_slave = performance_counter_0_control_slave_arb_winner[0] && cpu_3_data_master_requests_performance_counter_0_control_slave;

  //cpu_2/data_master assignment into master qualified-requests vector for performance_counter_0/control_slave, which is an e_assign
  assign performance_counter_0_control_slave_master_qreq_vector[1] = cpu_2_data_master_qualified_request_performance_counter_0_control_slave;

  //cpu_2/data_master grant performance_counter_0/control_slave, which is an e_assign
  assign cpu_2_data_master_granted_performance_counter_0_control_slave = performance_counter_0_control_slave_grant_vector[1];

  //cpu_2/data_master saved-grant performance_counter_0/control_slave, which is an e_assign
  assign cpu_2_data_master_saved_grant_performance_counter_0_control_slave = performance_counter_0_control_slave_arb_winner[1] && cpu_2_data_master_requests_performance_counter_0_control_slave;

  //cpu_1/data_master assignment into master qualified-requests vector for performance_counter_0/control_slave, which is an e_assign
  assign performance_counter_0_control_slave_master_qreq_vector[2] = cpu_1_data_master_qualified_request_performance_counter_0_control_slave;

  //cpu_1/data_master grant performance_counter_0/control_slave, which is an e_assign
  assign cpu_1_data_master_granted_performance_counter_0_control_slave = performance_counter_0_control_slave_grant_vector[2];

  //cpu_1/data_master saved-grant performance_counter_0/control_slave, which is an e_assign
  assign cpu_1_data_master_saved_grant_performance_counter_0_control_slave = performance_counter_0_control_slave_arb_winner[2] && cpu_1_data_master_requests_performance_counter_0_control_slave;

  //cpu_0/data_master assignment into master qualified-requests vector for performance_counter_0/control_slave, which is an e_assign
  assign performance_counter_0_control_slave_master_qreq_vector[3] = cpu_0_data_master_qualified_request_performance_counter_0_control_slave;

  //cpu_0/data_master grant performance_counter_0/control_slave, which is an e_assign
  assign cpu_0_data_master_granted_performance_counter_0_control_slave = performance_counter_0_control_slave_grant_vector[3];

  //cpu_0/data_master saved-grant performance_counter_0/control_slave, which is an e_assign
  assign cpu_0_data_master_saved_grant_performance_counter_0_control_slave = performance_counter_0_control_slave_arb_winner[3] && cpu_0_data_master_requests_performance_counter_0_control_slave;

  //performance_counter_0/control_slave chosen-master double-vector, which is an e_assign
  assign performance_counter_0_control_slave_chosen_master_double_vector = {performance_counter_0_control_slave_master_qreq_vector, performance_counter_0_control_slave_master_qreq_vector} & ({~performance_counter_0_control_slave_master_qreq_vector, ~performance_counter_0_control_slave_master_qreq_vector} + performance_counter_0_control_slave_arb_addend);

  //stable onehot encoding of arb winner
  assign performance_counter_0_control_slave_arb_winner = (performance_counter_0_control_slave_allow_new_arb_cycle & | performance_counter_0_control_slave_grant_vector) ? performance_counter_0_control_slave_grant_vector : performance_counter_0_control_slave_saved_chosen_master_vector;

  //saved performance_counter_0_control_slave_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          performance_counter_0_control_slave_saved_chosen_master_vector <= 0;
      else if (performance_counter_0_control_slave_allow_new_arb_cycle)
          performance_counter_0_control_slave_saved_chosen_master_vector <= |performance_counter_0_control_slave_grant_vector ? performance_counter_0_control_slave_grant_vector : performance_counter_0_control_slave_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign performance_counter_0_control_slave_grant_vector = {(performance_counter_0_control_slave_chosen_master_double_vector[3] | performance_counter_0_control_slave_chosen_master_double_vector[7]),
    (performance_counter_0_control_slave_chosen_master_double_vector[2] | performance_counter_0_control_slave_chosen_master_double_vector[6]),
    (performance_counter_0_control_slave_chosen_master_double_vector[1] | performance_counter_0_control_slave_chosen_master_double_vector[5]),
    (performance_counter_0_control_slave_chosen_master_double_vector[0] | performance_counter_0_control_slave_chosen_master_double_vector[4])};

  //performance_counter_0/control_slave chosen master rotated left, which is an e_assign
  assign performance_counter_0_control_slave_chosen_master_rot_left = (performance_counter_0_control_slave_arb_winner << 1) ? (performance_counter_0_control_slave_arb_winner << 1) : 1;

  //performance_counter_0/control_slave's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          performance_counter_0_control_slave_arb_addend <= 1;
      else if (|performance_counter_0_control_slave_grant_vector)
          performance_counter_0_control_slave_arb_addend <= performance_counter_0_control_slave_end_xfer? performance_counter_0_control_slave_chosen_master_rot_left : performance_counter_0_control_slave_grant_vector;
    end


  assign performance_counter_0_control_slave_begintransfer = performance_counter_0_control_slave_begins_xfer;
  //performance_counter_0_control_slave_reset_n assignment, which is an e_assign
  assign performance_counter_0_control_slave_reset_n = reset_n;

  //performance_counter_0_control_slave_firsttransfer first transaction, which is an e_assign
  assign performance_counter_0_control_slave_firsttransfer = performance_counter_0_control_slave_begins_xfer ? performance_counter_0_control_slave_unreg_firsttransfer : performance_counter_0_control_slave_reg_firsttransfer;

  //performance_counter_0_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign performance_counter_0_control_slave_unreg_firsttransfer = ~(performance_counter_0_control_slave_slavearbiterlockenable & performance_counter_0_control_slave_any_continuerequest);

  //performance_counter_0_control_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          performance_counter_0_control_slave_reg_firsttransfer <= 1'b1;
      else if (performance_counter_0_control_slave_begins_xfer)
          performance_counter_0_control_slave_reg_firsttransfer <= performance_counter_0_control_slave_unreg_firsttransfer;
    end


  //performance_counter_0_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign performance_counter_0_control_slave_beginbursttransfer_internal = performance_counter_0_control_slave_begins_xfer;

  //performance_counter_0_control_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign performance_counter_0_control_slave_arbitration_holdoff_internal = performance_counter_0_control_slave_begins_xfer & performance_counter_0_control_slave_firsttransfer;

  //performance_counter_0_control_slave_write assignment, which is an e_mux
  assign performance_counter_0_control_slave_write = (cpu_0_data_master_granted_performance_counter_0_control_slave & cpu_0_data_master_write) | (cpu_1_data_master_granted_performance_counter_0_control_slave & cpu_1_data_master_write) | (cpu_2_data_master_granted_performance_counter_0_control_slave & cpu_2_data_master_write) | (cpu_3_data_master_granted_performance_counter_0_control_slave & cpu_3_data_master_write);

  assign shifted_address_to_performance_counter_0_control_slave_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //performance_counter_0_control_slave_address mux, which is an e_mux
  assign performance_counter_0_control_slave_address = (cpu_0_data_master_granted_performance_counter_0_control_slave)? (shifted_address_to_performance_counter_0_control_slave_from_cpu_0_data_master >> 2) :
    (cpu_1_data_master_granted_performance_counter_0_control_slave)? (shifted_address_to_performance_counter_0_control_slave_from_cpu_1_data_master >> 2) :
    (cpu_2_data_master_granted_performance_counter_0_control_slave)? (shifted_address_to_performance_counter_0_control_slave_from_cpu_2_data_master >> 2) :
    (shifted_address_to_performance_counter_0_control_slave_from_cpu_3_data_master >> 2);

  assign shifted_address_to_performance_counter_0_control_slave_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_performance_counter_0_control_slave_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_performance_counter_0_control_slave_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  //d1_performance_counter_0_control_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_performance_counter_0_control_slave_end_xfer <= 1;
      else 
        d1_performance_counter_0_control_slave_end_xfer <= performance_counter_0_control_slave_end_xfer;
    end


  //performance_counter_0_control_slave_waits_for_read in a cycle, which is an e_mux
  assign performance_counter_0_control_slave_waits_for_read = performance_counter_0_control_slave_in_a_read_cycle & 0;

  //performance_counter_0_control_slave_in_a_read_cycle assignment, which is an e_assign
  assign performance_counter_0_control_slave_in_a_read_cycle = (cpu_0_data_master_granted_performance_counter_0_control_slave & cpu_0_data_master_read) | (cpu_1_data_master_granted_performance_counter_0_control_slave & cpu_1_data_master_read) | (cpu_2_data_master_granted_performance_counter_0_control_slave & cpu_2_data_master_read) | (cpu_3_data_master_granted_performance_counter_0_control_slave & cpu_3_data_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = performance_counter_0_control_slave_in_a_read_cycle;

  //performance_counter_0_control_slave_waits_for_write in a cycle, which is an e_mux
  assign performance_counter_0_control_slave_waits_for_write = performance_counter_0_control_slave_in_a_write_cycle & 0;

  //performance_counter_0_control_slave_in_a_write_cycle assignment, which is an e_assign
  assign performance_counter_0_control_slave_in_a_write_cycle = (cpu_0_data_master_granted_performance_counter_0_control_slave & cpu_0_data_master_write) | (cpu_1_data_master_granted_performance_counter_0_control_slave & cpu_1_data_master_write) | (cpu_2_data_master_granted_performance_counter_0_control_slave & cpu_2_data_master_write) | (cpu_3_data_master_granted_performance_counter_0_control_slave & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = performance_counter_0_control_slave_in_a_write_cycle;

  assign wait_for_performance_counter_0_control_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //performance_counter_0/control_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_performance_counter_0_control_slave + cpu_1_data_master_granted_performance_counter_0_control_slave + cpu_2_data_master_granted_performance_counter_0_control_slave + cpu_3_data_master_granted_performance_counter_0_control_slave > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_performance_counter_0_control_slave + cpu_1_data_master_saved_grant_performance_counter_0_control_slave + cpu_2_data_master_saved_grant_performance_counter_0_control_slave + cpu_3_data_master_saved_grant_performance_counter_0_control_slave > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_nios_system_clock_0_out_to_sdram_0_s1_module (
                                                                   // inputs:
                                                                    clear_fifo,
                                                                    clk,
                                                                    data_in,
                                                                    read,
                                                                    reset_n,
                                                                    sync_reset,
                                                                    write,

                                                                   // outputs:
                                                                    data_out,
                                                                    empty,
                                                                    fifo_contains_ones_n,
                                                                    full
                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_nios_system_clock_1_out_to_sdram_0_s1_module (
                                                                   // inputs:
                                                                    clear_fifo,
                                                                    clk,
                                                                    data_in,
                                                                    read,
                                                                    reset_n,
                                                                    sync_reset,
                                                                    write,

                                                                   // outputs:
                                                                    data_out,
                                                                    empty,
                                                                    fifo_contains_ones_n,
                                                                    full
                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_nios_system_clock_2_out_to_sdram_0_s1_module (
                                                                   // inputs:
                                                                    clear_fifo,
                                                                    clk,
                                                                    data_in,
                                                                    read,
                                                                    reset_n,
                                                                    sync_reset,
                                                                    write,

                                                                   // outputs:
                                                                    data_out,
                                                                    empty,
                                                                    fifo_contains_ones_n,
                                                                    full
                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_nios_system_clock_3_out_to_sdram_0_s1_module (
                                                                   // inputs:
                                                                    clear_fifo,
                                                                    clk,
                                                                    data_in,
                                                                    read,
                                                                    reset_n,
                                                                    sync_reset,
                                                                    write,

                                                                   // outputs:
                                                                    data_out,
                                                                    empty,
                                                                    fifo_contains_ones_n,
                                                                    full
                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_nios_system_clock_4_out_to_sdram_0_s1_module (
                                                                   // inputs:
                                                                    clear_fifo,
                                                                    clk,
                                                                    data_in,
                                                                    read,
                                                                    reset_n,
                                                                    sync_reset,
                                                                    write,

                                                                   // outputs:
                                                                    data_out,
                                                                    empty,
                                                                    fifo_contains_ones_n,
                                                                    full
                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_nios_system_clock_5_out_to_sdram_0_s1_module (
                                                                   // inputs:
                                                                    clear_fifo,
                                                                    clk,
                                                                    data_in,
                                                                    read,
                                                                    reset_n,
                                                                    sync_reset,
                                                                    write,

                                                                   // outputs:
                                                                    data_out,
                                                                    empty,
                                                                    fifo_contains_ones_n,
                                                                    full
                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_nios_system_clock_6_out_to_sdram_0_s1_module (
                                                                   // inputs:
                                                                    clear_fifo,
                                                                    clk,
                                                                    data_in,
                                                                    read,
                                                                    reset_n,
                                                                    sync_reset,
                                                                    write,

                                                                   // outputs:
                                                                    data_out,
                                                                    empty,
                                                                    fifo_contains_ones_n,
                                                                    full
                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_nios_system_clock_7_out_to_sdram_0_s1_module (
                                                                   // inputs:
                                                                    clear_fifo,
                                                                    clk,
                                                                    data_in,
                                                                    read,
                                                                    reset_n,
                                                                    sync_reset,
                                                                    write,

                                                                   // outputs:
                                                                    data_out,
                                                                    empty,
                                                                    fifo_contains_ones_n,
                                                                    full
                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sdram_0_s1_arbitrator (
                               // inputs:
                                clk,
                                nios_system_clock_0_out_address_to_slave,
                                nios_system_clock_0_out_byteenable,
                                nios_system_clock_0_out_read,
                                nios_system_clock_0_out_write,
                                nios_system_clock_0_out_writedata,
                                nios_system_clock_1_out_address_to_slave,
                                nios_system_clock_1_out_byteenable,
                                nios_system_clock_1_out_read,
                                nios_system_clock_1_out_write,
                                nios_system_clock_1_out_writedata,
                                nios_system_clock_2_out_address_to_slave,
                                nios_system_clock_2_out_byteenable,
                                nios_system_clock_2_out_read,
                                nios_system_clock_2_out_write,
                                nios_system_clock_2_out_writedata,
                                nios_system_clock_3_out_address_to_slave,
                                nios_system_clock_3_out_byteenable,
                                nios_system_clock_3_out_read,
                                nios_system_clock_3_out_write,
                                nios_system_clock_3_out_writedata,
                                nios_system_clock_4_out_address_to_slave,
                                nios_system_clock_4_out_byteenable,
                                nios_system_clock_4_out_read,
                                nios_system_clock_4_out_write,
                                nios_system_clock_4_out_writedata,
                                nios_system_clock_5_out_address_to_slave,
                                nios_system_clock_5_out_byteenable,
                                nios_system_clock_5_out_read,
                                nios_system_clock_5_out_write,
                                nios_system_clock_5_out_writedata,
                                nios_system_clock_6_out_address_to_slave,
                                nios_system_clock_6_out_byteenable,
                                nios_system_clock_6_out_read,
                                nios_system_clock_6_out_write,
                                nios_system_clock_6_out_writedata,
                                nios_system_clock_7_out_address_to_slave,
                                nios_system_clock_7_out_byteenable,
                                nios_system_clock_7_out_read,
                                nios_system_clock_7_out_write,
                                nios_system_clock_7_out_writedata,
                                reset_n,
                                sdram_0_s1_readdata,
                                sdram_0_s1_readdatavalid,
                                sdram_0_s1_waitrequest,

                               // outputs:
                                d1_sdram_0_s1_end_xfer,
                                nios_system_clock_0_out_granted_sdram_0_s1,
                                nios_system_clock_0_out_qualified_request_sdram_0_s1,
                                nios_system_clock_0_out_read_data_valid_sdram_0_s1,
                                nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register,
                                nios_system_clock_0_out_requests_sdram_0_s1,
                                nios_system_clock_1_out_granted_sdram_0_s1,
                                nios_system_clock_1_out_qualified_request_sdram_0_s1,
                                nios_system_clock_1_out_read_data_valid_sdram_0_s1,
                                nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register,
                                nios_system_clock_1_out_requests_sdram_0_s1,
                                nios_system_clock_2_out_granted_sdram_0_s1,
                                nios_system_clock_2_out_qualified_request_sdram_0_s1,
                                nios_system_clock_2_out_read_data_valid_sdram_0_s1,
                                nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register,
                                nios_system_clock_2_out_requests_sdram_0_s1,
                                nios_system_clock_3_out_granted_sdram_0_s1,
                                nios_system_clock_3_out_qualified_request_sdram_0_s1,
                                nios_system_clock_3_out_read_data_valid_sdram_0_s1,
                                nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register,
                                nios_system_clock_3_out_requests_sdram_0_s1,
                                nios_system_clock_4_out_granted_sdram_0_s1,
                                nios_system_clock_4_out_qualified_request_sdram_0_s1,
                                nios_system_clock_4_out_read_data_valid_sdram_0_s1,
                                nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register,
                                nios_system_clock_4_out_requests_sdram_0_s1,
                                nios_system_clock_5_out_granted_sdram_0_s1,
                                nios_system_clock_5_out_qualified_request_sdram_0_s1,
                                nios_system_clock_5_out_read_data_valid_sdram_0_s1,
                                nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register,
                                nios_system_clock_5_out_requests_sdram_0_s1,
                                nios_system_clock_6_out_granted_sdram_0_s1,
                                nios_system_clock_6_out_qualified_request_sdram_0_s1,
                                nios_system_clock_6_out_read_data_valid_sdram_0_s1,
                                nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register,
                                nios_system_clock_6_out_requests_sdram_0_s1,
                                nios_system_clock_7_out_granted_sdram_0_s1,
                                nios_system_clock_7_out_qualified_request_sdram_0_s1,
                                nios_system_clock_7_out_read_data_valid_sdram_0_s1,
                                nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register,
                                nios_system_clock_7_out_requests_sdram_0_s1,
                                sdram_0_s1_address,
                                sdram_0_s1_byteenable_n,
                                sdram_0_s1_chipselect,
                                sdram_0_s1_read_n,
                                sdram_0_s1_readdata_from_sa,
                                sdram_0_s1_reset_n,
                                sdram_0_s1_waitrequest_from_sa,
                                sdram_0_s1_write_n,
                                sdram_0_s1_writedata
                             )
;

  output           d1_sdram_0_s1_end_xfer;
  output           nios_system_clock_0_out_granted_sdram_0_s1;
  output           nios_system_clock_0_out_qualified_request_sdram_0_s1;
  output           nios_system_clock_0_out_read_data_valid_sdram_0_s1;
  output           nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register;
  output           nios_system_clock_0_out_requests_sdram_0_s1;
  output           nios_system_clock_1_out_granted_sdram_0_s1;
  output           nios_system_clock_1_out_qualified_request_sdram_0_s1;
  output           nios_system_clock_1_out_read_data_valid_sdram_0_s1;
  output           nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register;
  output           nios_system_clock_1_out_requests_sdram_0_s1;
  output           nios_system_clock_2_out_granted_sdram_0_s1;
  output           nios_system_clock_2_out_qualified_request_sdram_0_s1;
  output           nios_system_clock_2_out_read_data_valid_sdram_0_s1;
  output           nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register;
  output           nios_system_clock_2_out_requests_sdram_0_s1;
  output           nios_system_clock_3_out_granted_sdram_0_s1;
  output           nios_system_clock_3_out_qualified_request_sdram_0_s1;
  output           nios_system_clock_3_out_read_data_valid_sdram_0_s1;
  output           nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register;
  output           nios_system_clock_3_out_requests_sdram_0_s1;
  output           nios_system_clock_4_out_granted_sdram_0_s1;
  output           nios_system_clock_4_out_qualified_request_sdram_0_s1;
  output           nios_system_clock_4_out_read_data_valid_sdram_0_s1;
  output           nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register;
  output           nios_system_clock_4_out_requests_sdram_0_s1;
  output           nios_system_clock_5_out_granted_sdram_0_s1;
  output           nios_system_clock_5_out_qualified_request_sdram_0_s1;
  output           nios_system_clock_5_out_read_data_valid_sdram_0_s1;
  output           nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register;
  output           nios_system_clock_5_out_requests_sdram_0_s1;
  output           nios_system_clock_6_out_granted_sdram_0_s1;
  output           nios_system_clock_6_out_qualified_request_sdram_0_s1;
  output           nios_system_clock_6_out_read_data_valid_sdram_0_s1;
  output           nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register;
  output           nios_system_clock_6_out_requests_sdram_0_s1;
  output           nios_system_clock_7_out_granted_sdram_0_s1;
  output           nios_system_clock_7_out_qualified_request_sdram_0_s1;
  output           nios_system_clock_7_out_read_data_valid_sdram_0_s1;
  output           nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register;
  output           nios_system_clock_7_out_requests_sdram_0_s1;
  output  [ 21: 0] sdram_0_s1_address;
  output  [  1: 0] sdram_0_s1_byteenable_n;
  output           sdram_0_s1_chipselect;
  output           sdram_0_s1_read_n;
  output  [ 15: 0] sdram_0_s1_readdata_from_sa;
  output           sdram_0_s1_reset_n;
  output           sdram_0_s1_waitrequest_from_sa;
  output           sdram_0_s1_write_n;
  output  [ 15: 0] sdram_0_s1_writedata;
  input            clk;
  input   [ 22: 0] nios_system_clock_0_out_address_to_slave;
  input   [  1: 0] nios_system_clock_0_out_byteenable;
  input            nios_system_clock_0_out_read;
  input            nios_system_clock_0_out_write;
  input   [ 15: 0] nios_system_clock_0_out_writedata;
  input   [ 22: 0] nios_system_clock_1_out_address_to_slave;
  input   [  1: 0] nios_system_clock_1_out_byteenable;
  input            nios_system_clock_1_out_read;
  input            nios_system_clock_1_out_write;
  input   [ 15: 0] nios_system_clock_1_out_writedata;
  input   [ 22: 0] nios_system_clock_2_out_address_to_slave;
  input   [  1: 0] nios_system_clock_2_out_byteenable;
  input            nios_system_clock_2_out_read;
  input            nios_system_clock_2_out_write;
  input   [ 15: 0] nios_system_clock_2_out_writedata;
  input   [ 22: 0] nios_system_clock_3_out_address_to_slave;
  input   [  1: 0] nios_system_clock_3_out_byteenable;
  input            nios_system_clock_3_out_read;
  input            nios_system_clock_3_out_write;
  input   [ 15: 0] nios_system_clock_3_out_writedata;
  input   [ 22: 0] nios_system_clock_4_out_address_to_slave;
  input   [  1: 0] nios_system_clock_4_out_byteenable;
  input            nios_system_clock_4_out_read;
  input            nios_system_clock_4_out_write;
  input   [ 15: 0] nios_system_clock_4_out_writedata;
  input   [ 22: 0] nios_system_clock_5_out_address_to_slave;
  input   [  1: 0] nios_system_clock_5_out_byteenable;
  input            nios_system_clock_5_out_read;
  input            nios_system_clock_5_out_write;
  input   [ 15: 0] nios_system_clock_5_out_writedata;
  input   [ 22: 0] nios_system_clock_6_out_address_to_slave;
  input   [  1: 0] nios_system_clock_6_out_byteenable;
  input            nios_system_clock_6_out_read;
  input            nios_system_clock_6_out_write;
  input   [ 15: 0] nios_system_clock_6_out_writedata;
  input   [ 22: 0] nios_system_clock_7_out_address_to_slave;
  input   [  1: 0] nios_system_clock_7_out_byteenable;
  input            nios_system_clock_7_out_read;
  input            nios_system_clock_7_out_write;
  input   [ 15: 0] nios_system_clock_7_out_writedata;
  input            reset_n;
  input   [ 15: 0] sdram_0_s1_readdata;
  input            sdram_0_s1_readdatavalid;
  input            sdram_0_s1_waitrequest;

  reg              d1_reasons_to_wait;
  reg              d1_sdram_0_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sdram_0_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_nios_system_clock_0_out_granted_slave_sdram_0_s1;
  reg              last_cycle_nios_system_clock_1_out_granted_slave_sdram_0_s1;
  reg              last_cycle_nios_system_clock_2_out_granted_slave_sdram_0_s1;
  reg              last_cycle_nios_system_clock_3_out_granted_slave_sdram_0_s1;
  reg              last_cycle_nios_system_clock_4_out_granted_slave_sdram_0_s1;
  reg              last_cycle_nios_system_clock_5_out_granted_slave_sdram_0_s1;
  reg              last_cycle_nios_system_clock_6_out_granted_slave_sdram_0_s1;
  reg              last_cycle_nios_system_clock_7_out_granted_slave_sdram_0_s1;
  wire             nios_system_clock_0_out_arbiterlock;
  wire             nios_system_clock_0_out_arbiterlock2;
  wire             nios_system_clock_0_out_continuerequest;
  wire             nios_system_clock_0_out_granted_sdram_0_s1;
  wire             nios_system_clock_0_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_0_out_rdv_fifo_empty_sdram_0_s1;
  wire             nios_system_clock_0_out_rdv_fifo_output_from_sdram_0_s1;
  wire             nios_system_clock_0_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register;
  wire             nios_system_clock_0_out_requests_sdram_0_s1;
  wire             nios_system_clock_0_out_saved_grant_sdram_0_s1;
  wire             nios_system_clock_1_out_arbiterlock;
  wire             nios_system_clock_1_out_arbiterlock2;
  wire             nios_system_clock_1_out_continuerequest;
  wire             nios_system_clock_1_out_granted_sdram_0_s1;
  wire             nios_system_clock_1_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_1_out_rdv_fifo_empty_sdram_0_s1;
  wire             nios_system_clock_1_out_rdv_fifo_output_from_sdram_0_s1;
  wire             nios_system_clock_1_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register;
  wire             nios_system_clock_1_out_requests_sdram_0_s1;
  wire             nios_system_clock_1_out_saved_grant_sdram_0_s1;
  wire             nios_system_clock_2_out_arbiterlock;
  wire             nios_system_clock_2_out_arbiterlock2;
  wire             nios_system_clock_2_out_continuerequest;
  wire             nios_system_clock_2_out_granted_sdram_0_s1;
  wire             nios_system_clock_2_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_2_out_rdv_fifo_empty_sdram_0_s1;
  wire             nios_system_clock_2_out_rdv_fifo_output_from_sdram_0_s1;
  wire             nios_system_clock_2_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register;
  wire             nios_system_clock_2_out_requests_sdram_0_s1;
  wire             nios_system_clock_2_out_saved_grant_sdram_0_s1;
  wire             nios_system_clock_3_out_arbiterlock;
  wire             nios_system_clock_3_out_arbiterlock2;
  wire             nios_system_clock_3_out_continuerequest;
  wire             nios_system_clock_3_out_granted_sdram_0_s1;
  wire             nios_system_clock_3_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_3_out_rdv_fifo_empty_sdram_0_s1;
  wire             nios_system_clock_3_out_rdv_fifo_output_from_sdram_0_s1;
  wire             nios_system_clock_3_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register;
  wire             nios_system_clock_3_out_requests_sdram_0_s1;
  wire             nios_system_clock_3_out_saved_grant_sdram_0_s1;
  wire             nios_system_clock_4_out_arbiterlock;
  wire             nios_system_clock_4_out_arbiterlock2;
  wire             nios_system_clock_4_out_continuerequest;
  wire             nios_system_clock_4_out_granted_sdram_0_s1;
  wire             nios_system_clock_4_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_4_out_rdv_fifo_empty_sdram_0_s1;
  wire             nios_system_clock_4_out_rdv_fifo_output_from_sdram_0_s1;
  wire             nios_system_clock_4_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register;
  wire             nios_system_clock_4_out_requests_sdram_0_s1;
  wire             nios_system_clock_4_out_saved_grant_sdram_0_s1;
  wire             nios_system_clock_5_out_arbiterlock;
  wire             nios_system_clock_5_out_arbiterlock2;
  wire             nios_system_clock_5_out_continuerequest;
  wire             nios_system_clock_5_out_granted_sdram_0_s1;
  wire             nios_system_clock_5_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_5_out_rdv_fifo_empty_sdram_0_s1;
  wire             nios_system_clock_5_out_rdv_fifo_output_from_sdram_0_s1;
  wire             nios_system_clock_5_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register;
  wire             nios_system_clock_5_out_requests_sdram_0_s1;
  wire             nios_system_clock_5_out_saved_grant_sdram_0_s1;
  wire             nios_system_clock_6_out_arbiterlock;
  wire             nios_system_clock_6_out_arbiterlock2;
  wire             nios_system_clock_6_out_continuerequest;
  wire             nios_system_clock_6_out_granted_sdram_0_s1;
  wire             nios_system_clock_6_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_6_out_rdv_fifo_empty_sdram_0_s1;
  wire             nios_system_clock_6_out_rdv_fifo_output_from_sdram_0_s1;
  wire             nios_system_clock_6_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register;
  wire             nios_system_clock_6_out_requests_sdram_0_s1;
  wire             nios_system_clock_6_out_saved_grant_sdram_0_s1;
  wire             nios_system_clock_7_out_arbiterlock;
  wire             nios_system_clock_7_out_arbiterlock2;
  wire             nios_system_clock_7_out_continuerequest;
  wire             nios_system_clock_7_out_granted_sdram_0_s1;
  wire             nios_system_clock_7_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_7_out_rdv_fifo_empty_sdram_0_s1;
  wire             nios_system_clock_7_out_rdv_fifo_output_from_sdram_0_s1;
  wire             nios_system_clock_7_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register;
  wire             nios_system_clock_7_out_requests_sdram_0_s1;
  wire             nios_system_clock_7_out_saved_grant_sdram_0_s1;
  wire    [ 21: 0] sdram_0_s1_address;
  wire             sdram_0_s1_allgrants;
  wire             sdram_0_s1_allow_new_arb_cycle;
  wire             sdram_0_s1_any_bursting_master_saved_grant;
  wire             sdram_0_s1_any_continuerequest;
  reg     [  7: 0] sdram_0_s1_arb_addend;
  wire             sdram_0_s1_arb_counter_enable;
  reg              sdram_0_s1_arb_share_counter;
  wire             sdram_0_s1_arb_share_counter_next_value;
  wire             sdram_0_s1_arb_share_set_values;
  wire    [  7: 0] sdram_0_s1_arb_winner;
  wire             sdram_0_s1_arbitration_holdoff_internal;
  wire             sdram_0_s1_beginbursttransfer_internal;
  wire             sdram_0_s1_begins_xfer;
  wire    [  1: 0] sdram_0_s1_byteenable_n;
  wire             sdram_0_s1_chipselect;
  wire    [ 15: 0] sdram_0_s1_chosen_master_double_vector;
  wire    [  7: 0] sdram_0_s1_chosen_master_rot_left;
  wire             sdram_0_s1_end_xfer;
  wire             sdram_0_s1_firsttransfer;
  wire    [  7: 0] sdram_0_s1_grant_vector;
  wire             sdram_0_s1_in_a_read_cycle;
  wire             sdram_0_s1_in_a_write_cycle;
  wire    [  7: 0] sdram_0_s1_master_qreq_vector;
  wire             sdram_0_s1_move_on_to_next_transaction;
  wire             sdram_0_s1_non_bursting_master_requests;
  wire             sdram_0_s1_read_n;
  wire    [ 15: 0] sdram_0_s1_readdata_from_sa;
  wire             sdram_0_s1_readdatavalid_from_sa;
  reg              sdram_0_s1_reg_firsttransfer;
  wire             sdram_0_s1_reset_n;
  reg     [  7: 0] sdram_0_s1_saved_chosen_master_vector;
  reg              sdram_0_s1_slavearbiterlockenable;
  wire             sdram_0_s1_slavearbiterlockenable2;
  wire             sdram_0_s1_unreg_firsttransfer;
  wire             sdram_0_s1_waitrequest_from_sa;
  wire             sdram_0_s1_waits_for_read;
  wire             sdram_0_s1_waits_for_write;
  wire             sdram_0_s1_write_n;
  wire    [ 15: 0] sdram_0_s1_writedata;
  wire    [ 22: 0] shifted_address_to_sdram_0_s1_from_nios_system_clock_0_out;
  wire    [ 22: 0] shifted_address_to_sdram_0_s1_from_nios_system_clock_1_out;
  wire    [ 22: 0] shifted_address_to_sdram_0_s1_from_nios_system_clock_2_out;
  wire    [ 22: 0] shifted_address_to_sdram_0_s1_from_nios_system_clock_3_out;
  wire    [ 22: 0] shifted_address_to_sdram_0_s1_from_nios_system_clock_4_out;
  wire    [ 22: 0] shifted_address_to_sdram_0_s1_from_nios_system_clock_5_out;
  wire    [ 22: 0] shifted_address_to_sdram_0_s1_from_nios_system_clock_6_out;
  wire    [ 22: 0] shifted_address_to_sdram_0_s1_from_nios_system_clock_7_out;
  wire             wait_for_sdram_0_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sdram_0_s1_end_xfer;
    end


  assign sdram_0_s1_begins_xfer = ~d1_reasons_to_wait & ((nios_system_clock_0_out_qualified_request_sdram_0_s1 | nios_system_clock_1_out_qualified_request_sdram_0_s1 | nios_system_clock_2_out_qualified_request_sdram_0_s1 | nios_system_clock_3_out_qualified_request_sdram_0_s1 | nios_system_clock_4_out_qualified_request_sdram_0_s1 | nios_system_clock_5_out_qualified_request_sdram_0_s1 | nios_system_clock_6_out_qualified_request_sdram_0_s1 | nios_system_clock_7_out_qualified_request_sdram_0_s1));
  //assign sdram_0_s1_readdata_from_sa = sdram_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_0_s1_readdata_from_sa = sdram_0_s1_readdata;

  assign nios_system_clock_0_out_requests_sdram_0_s1 = (1) & (nios_system_clock_0_out_read | nios_system_clock_0_out_write);
  //assign sdram_0_s1_waitrequest_from_sa = sdram_0_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_0_s1_waitrequest_from_sa = sdram_0_s1_waitrequest;

  //assign sdram_0_s1_readdatavalid_from_sa = sdram_0_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_0_s1_readdatavalid_from_sa = sdram_0_s1_readdatavalid;

  //sdram_0_s1_arb_share_counter set values, which is an e_mux
  assign sdram_0_s1_arb_share_set_values = 1;

  //sdram_0_s1_non_bursting_master_requests mux, which is an e_mux
  assign sdram_0_s1_non_bursting_master_requests = nios_system_clock_0_out_requests_sdram_0_s1 |
    nios_system_clock_1_out_requests_sdram_0_s1 |
    nios_system_clock_2_out_requests_sdram_0_s1 |
    nios_system_clock_3_out_requests_sdram_0_s1 |
    nios_system_clock_4_out_requests_sdram_0_s1 |
    nios_system_clock_5_out_requests_sdram_0_s1 |
    nios_system_clock_6_out_requests_sdram_0_s1 |
    nios_system_clock_7_out_requests_sdram_0_s1 |
    nios_system_clock_0_out_requests_sdram_0_s1 |
    nios_system_clock_1_out_requests_sdram_0_s1 |
    nios_system_clock_2_out_requests_sdram_0_s1 |
    nios_system_clock_3_out_requests_sdram_0_s1 |
    nios_system_clock_4_out_requests_sdram_0_s1 |
    nios_system_clock_5_out_requests_sdram_0_s1 |
    nios_system_clock_6_out_requests_sdram_0_s1 |
    nios_system_clock_7_out_requests_sdram_0_s1 |
    nios_system_clock_0_out_requests_sdram_0_s1 |
    nios_system_clock_1_out_requests_sdram_0_s1 |
    nios_system_clock_2_out_requests_sdram_0_s1 |
    nios_system_clock_3_out_requests_sdram_0_s1 |
    nios_system_clock_4_out_requests_sdram_0_s1 |
    nios_system_clock_5_out_requests_sdram_0_s1 |
    nios_system_clock_6_out_requests_sdram_0_s1 |
    nios_system_clock_7_out_requests_sdram_0_s1 |
    nios_system_clock_0_out_requests_sdram_0_s1 |
    nios_system_clock_1_out_requests_sdram_0_s1 |
    nios_system_clock_2_out_requests_sdram_0_s1 |
    nios_system_clock_3_out_requests_sdram_0_s1 |
    nios_system_clock_4_out_requests_sdram_0_s1 |
    nios_system_clock_5_out_requests_sdram_0_s1 |
    nios_system_clock_6_out_requests_sdram_0_s1 |
    nios_system_clock_7_out_requests_sdram_0_s1 |
    nios_system_clock_0_out_requests_sdram_0_s1 |
    nios_system_clock_1_out_requests_sdram_0_s1 |
    nios_system_clock_2_out_requests_sdram_0_s1 |
    nios_system_clock_3_out_requests_sdram_0_s1 |
    nios_system_clock_4_out_requests_sdram_0_s1 |
    nios_system_clock_5_out_requests_sdram_0_s1 |
    nios_system_clock_6_out_requests_sdram_0_s1 |
    nios_system_clock_7_out_requests_sdram_0_s1 |
    nios_system_clock_0_out_requests_sdram_0_s1 |
    nios_system_clock_1_out_requests_sdram_0_s1 |
    nios_system_clock_2_out_requests_sdram_0_s1 |
    nios_system_clock_3_out_requests_sdram_0_s1 |
    nios_system_clock_4_out_requests_sdram_0_s1 |
    nios_system_clock_5_out_requests_sdram_0_s1 |
    nios_system_clock_6_out_requests_sdram_0_s1 |
    nios_system_clock_7_out_requests_sdram_0_s1 |
    nios_system_clock_0_out_requests_sdram_0_s1 |
    nios_system_clock_1_out_requests_sdram_0_s1 |
    nios_system_clock_2_out_requests_sdram_0_s1 |
    nios_system_clock_3_out_requests_sdram_0_s1 |
    nios_system_clock_4_out_requests_sdram_0_s1 |
    nios_system_clock_5_out_requests_sdram_0_s1 |
    nios_system_clock_6_out_requests_sdram_0_s1 |
    nios_system_clock_7_out_requests_sdram_0_s1 |
    nios_system_clock_0_out_requests_sdram_0_s1 |
    nios_system_clock_1_out_requests_sdram_0_s1 |
    nios_system_clock_2_out_requests_sdram_0_s1 |
    nios_system_clock_3_out_requests_sdram_0_s1 |
    nios_system_clock_4_out_requests_sdram_0_s1 |
    nios_system_clock_5_out_requests_sdram_0_s1 |
    nios_system_clock_6_out_requests_sdram_0_s1 |
    nios_system_clock_7_out_requests_sdram_0_s1;

  //sdram_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign sdram_0_s1_any_bursting_master_saved_grant = 0;

  //sdram_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign sdram_0_s1_arb_share_counter_next_value = sdram_0_s1_firsttransfer ? (sdram_0_s1_arb_share_set_values - 1) : |sdram_0_s1_arb_share_counter ? (sdram_0_s1_arb_share_counter - 1) : 0;

  //sdram_0_s1_allgrants all slave grants, which is an e_mux
  assign sdram_0_s1_allgrants = (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector);

  //sdram_0_s1_end_xfer assignment, which is an e_assign
  assign sdram_0_s1_end_xfer = ~(sdram_0_s1_waits_for_read | sdram_0_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_sdram_0_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sdram_0_s1 = sdram_0_s1_end_xfer & (~sdram_0_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sdram_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign sdram_0_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_sdram_0_s1 & sdram_0_s1_allgrants) | (end_xfer_arb_share_counter_term_sdram_0_s1 & ~sdram_0_s1_non_bursting_master_requests);

  //sdram_0_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_0_s1_arb_share_counter <= 0;
      else if (sdram_0_s1_arb_counter_enable)
          sdram_0_s1_arb_share_counter <= sdram_0_s1_arb_share_counter_next_value;
    end


  //sdram_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_0_s1_slavearbiterlockenable <= 0;
      else if ((|sdram_0_s1_master_qreq_vector & end_xfer_arb_share_counter_term_sdram_0_s1) | (end_xfer_arb_share_counter_term_sdram_0_s1 & ~sdram_0_s1_non_bursting_master_requests))
          sdram_0_s1_slavearbiterlockenable <= |sdram_0_s1_arb_share_counter_next_value;
    end


  //nios_system_clock_0/out sdram_0/s1 arbiterlock, which is an e_assign
  assign nios_system_clock_0_out_arbiterlock = sdram_0_s1_slavearbiterlockenable & nios_system_clock_0_out_continuerequest;

  //sdram_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sdram_0_s1_slavearbiterlockenable2 = |sdram_0_s1_arb_share_counter_next_value;

  //nios_system_clock_0/out sdram_0/s1 arbiterlock2, which is an e_assign
  assign nios_system_clock_0_out_arbiterlock2 = sdram_0_s1_slavearbiterlockenable2 & nios_system_clock_0_out_continuerequest;

  //nios_system_clock_1/out sdram_0/s1 arbiterlock, which is an e_assign
  assign nios_system_clock_1_out_arbiterlock = sdram_0_s1_slavearbiterlockenable & nios_system_clock_1_out_continuerequest;

  //nios_system_clock_1/out sdram_0/s1 arbiterlock2, which is an e_assign
  assign nios_system_clock_1_out_arbiterlock2 = sdram_0_s1_slavearbiterlockenable2 & nios_system_clock_1_out_continuerequest;

  //nios_system_clock_1/out granted sdram_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_1_out_granted_slave_sdram_0_s1 <= 0;
      else 
        last_cycle_nios_system_clock_1_out_granted_slave_sdram_0_s1 <= nios_system_clock_1_out_saved_grant_sdram_0_s1 ? 1 : (sdram_0_s1_arbitration_holdoff_internal | ~nios_system_clock_1_out_requests_sdram_0_s1) ? 0 : last_cycle_nios_system_clock_1_out_granted_slave_sdram_0_s1;
    end


  //nios_system_clock_1_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_1_out_continuerequest = (last_cycle_nios_system_clock_1_out_granted_slave_sdram_0_s1 & nios_system_clock_1_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_1_out_granted_slave_sdram_0_s1 & nios_system_clock_1_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_1_out_granted_slave_sdram_0_s1 & nios_system_clock_1_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_1_out_granted_slave_sdram_0_s1 & nios_system_clock_1_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_1_out_granted_slave_sdram_0_s1 & nios_system_clock_1_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_1_out_granted_slave_sdram_0_s1 & nios_system_clock_1_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_1_out_granted_slave_sdram_0_s1 & nios_system_clock_1_out_requests_sdram_0_s1);

  //sdram_0_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign sdram_0_s1_any_continuerequest = nios_system_clock_1_out_continuerequest |
    nios_system_clock_2_out_continuerequest |
    nios_system_clock_3_out_continuerequest |
    nios_system_clock_4_out_continuerequest |
    nios_system_clock_5_out_continuerequest |
    nios_system_clock_6_out_continuerequest |
    nios_system_clock_7_out_continuerequest |
    nios_system_clock_0_out_continuerequest |
    nios_system_clock_2_out_continuerequest |
    nios_system_clock_3_out_continuerequest |
    nios_system_clock_4_out_continuerequest |
    nios_system_clock_5_out_continuerequest |
    nios_system_clock_6_out_continuerequest |
    nios_system_clock_7_out_continuerequest |
    nios_system_clock_0_out_continuerequest |
    nios_system_clock_1_out_continuerequest |
    nios_system_clock_3_out_continuerequest |
    nios_system_clock_4_out_continuerequest |
    nios_system_clock_5_out_continuerequest |
    nios_system_clock_6_out_continuerequest |
    nios_system_clock_7_out_continuerequest |
    nios_system_clock_0_out_continuerequest |
    nios_system_clock_1_out_continuerequest |
    nios_system_clock_2_out_continuerequest |
    nios_system_clock_4_out_continuerequest |
    nios_system_clock_5_out_continuerequest |
    nios_system_clock_6_out_continuerequest |
    nios_system_clock_7_out_continuerequest |
    nios_system_clock_0_out_continuerequest |
    nios_system_clock_1_out_continuerequest |
    nios_system_clock_2_out_continuerequest |
    nios_system_clock_3_out_continuerequest |
    nios_system_clock_5_out_continuerequest |
    nios_system_clock_6_out_continuerequest |
    nios_system_clock_7_out_continuerequest |
    nios_system_clock_0_out_continuerequest |
    nios_system_clock_1_out_continuerequest |
    nios_system_clock_2_out_continuerequest |
    nios_system_clock_3_out_continuerequest |
    nios_system_clock_4_out_continuerequest |
    nios_system_clock_6_out_continuerequest |
    nios_system_clock_7_out_continuerequest |
    nios_system_clock_0_out_continuerequest |
    nios_system_clock_1_out_continuerequest |
    nios_system_clock_2_out_continuerequest |
    nios_system_clock_3_out_continuerequest |
    nios_system_clock_4_out_continuerequest |
    nios_system_clock_5_out_continuerequest |
    nios_system_clock_7_out_continuerequest |
    nios_system_clock_0_out_continuerequest |
    nios_system_clock_1_out_continuerequest |
    nios_system_clock_2_out_continuerequest |
    nios_system_clock_3_out_continuerequest |
    nios_system_clock_4_out_continuerequest |
    nios_system_clock_5_out_continuerequest |
    nios_system_clock_6_out_continuerequest;

  //nios_system_clock_2/out sdram_0/s1 arbiterlock, which is an e_assign
  assign nios_system_clock_2_out_arbiterlock = sdram_0_s1_slavearbiterlockenable & nios_system_clock_2_out_continuerequest;

  //nios_system_clock_2/out sdram_0/s1 arbiterlock2, which is an e_assign
  assign nios_system_clock_2_out_arbiterlock2 = sdram_0_s1_slavearbiterlockenable2 & nios_system_clock_2_out_continuerequest;

  //nios_system_clock_2/out granted sdram_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_2_out_granted_slave_sdram_0_s1 <= 0;
      else 
        last_cycle_nios_system_clock_2_out_granted_slave_sdram_0_s1 <= nios_system_clock_2_out_saved_grant_sdram_0_s1 ? 1 : (sdram_0_s1_arbitration_holdoff_internal | ~nios_system_clock_2_out_requests_sdram_0_s1) ? 0 : last_cycle_nios_system_clock_2_out_granted_slave_sdram_0_s1;
    end


  //nios_system_clock_2_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_2_out_continuerequest = (last_cycle_nios_system_clock_2_out_granted_slave_sdram_0_s1 & nios_system_clock_2_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_2_out_granted_slave_sdram_0_s1 & nios_system_clock_2_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_2_out_granted_slave_sdram_0_s1 & nios_system_clock_2_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_2_out_granted_slave_sdram_0_s1 & nios_system_clock_2_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_2_out_granted_slave_sdram_0_s1 & nios_system_clock_2_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_2_out_granted_slave_sdram_0_s1 & nios_system_clock_2_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_2_out_granted_slave_sdram_0_s1 & nios_system_clock_2_out_requests_sdram_0_s1);

  //nios_system_clock_3/out sdram_0/s1 arbiterlock, which is an e_assign
  assign nios_system_clock_3_out_arbiterlock = sdram_0_s1_slavearbiterlockenable & nios_system_clock_3_out_continuerequest;

  //nios_system_clock_3/out sdram_0/s1 arbiterlock2, which is an e_assign
  assign nios_system_clock_3_out_arbiterlock2 = sdram_0_s1_slavearbiterlockenable2 & nios_system_clock_3_out_continuerequest;

  //nios_system_clock_3/out granted sdram_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_3_out_granted_slave_sdram_0_s1 <= 0;
      else 
        last_cycle_nios_system_clock_3_out_granted_slave_sdram_0_s1 <= nios_system_clock_3_out_saved_grant_sdram_0_s1 ? 1 : (sdram_0_s1_arbitration_holdoff_internal | ~nios_system_clock_3_out_requests_sdram_0_s1) ? 0 : last_cycle_nios_system_clock_3_out_granted_slave_sdram_0_s1;
    end


  //nios_system_clock_3_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_3_out_continuerequest = (last_cycle_nios_system_clock_3_out_granted_slave_sdram_0_s1 & nios_system_clock_3_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_3_out_granted_slave_sdram_0_s1 & nios_system_clock_3_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_3_out_granted_slave_sdram_0_s1 & nios_system_clock_3_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_3_out_granted_slave_sdram_0_s1 & nios_system_clock_3_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_3_out_granted_slave_sdram_0_s1 & nios_system_clock_3_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_3_out_granted_slave_sdram_0_s1 & nios_system_clock_3_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_3_out_granted_slave_sdram_0_s1 & nios_system_clock_3_out_requests_sdram_0_s1);

  //nios_system_clock_4/out sdram_0/s1 arbiterlock, which is an e_assign
  assign nios_system_clock_4_out_arbiterlock = sdram_0_s1_slavearbiterlockenable & nios_system_clock_4_out_continuerequest;

  //nios_system_clock_4/out sdram_0/s1 arbiterlock2, which is an e_assign
  assign nios_system_clock_4_out_arbiterlock2 = sdram_0_s1_slavearbiterlockenable2 & nios_system_clock_4_out_continuerequest;

  //nios_system_clock_4/out granted sdram_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_4_out_granted_slave_sdram_0_s1 <= 0;
      else 
        last_cycle_nios_system_clock_4_out_granted_slave_sdram_0_s1 <= nios_system_clock_4_out_saved_grant_sdram_0_s1 ? 1 : (sdram_0_s1_arbitration_holdoff_internal | ~nios_system_clock_4_out_requests_sdram_0_s1) ? 0 : last_cycle_nios_system_clock_4_out_granted_slave_sdram_0_s1;
    end


  //nios_system_clock_4_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_4_out_continuerequest = (last_cycle_nios_system_clock_4_out_granted_slave_sdram_0_s1 & nios_system_clock_4_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_4_out_granted_slave_sdram_0_s1 & nios_system_clock_4_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_4_out_granted_slave_sdram_0_s1 & nios_system_clock_4_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_4_out_granted_slave_sdram_0_s1 & nios_system_clock_4_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_4_out_granted_slave_sdram_0_s1 & nios_system_clock_4_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_4_out_granted_slave_sdram_0_s1 & nios_system_clock_4_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_4_out_granted_slave_sdram_0_s1 & nios_system_clock_4_out_requests_sdram_0_s1);

  //nios_system_clock_5/out sdram_0/s1 arbiterlock, which is an e_assign
  assign nios_system_clock_5_out_arbiterlock = sdram_0_s1_slavearbiterlockenable & nios_system_clock_5_out_continuerequest;

  //nios_system_clock_5/out sdram_0/s1 arbiterlock2, which is an e_assign
  assign nios_system_clock_5_out_arbiterlock2 = sdram_0_s1_slavearbiterlockenable2 & nios_system_clock_5_out_continuerequest;

  //nios_system_clock_5/out granted sdram_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_5_out_granted_slave_sdram_0_s1 <= 0;
      else 
        last_cycle_nios_system_clock_5_out_granted_slave_sdram_0_s1 <= nios_system_clock_5_out_saved_grant_sdram_0_s1 ? 1 : (sdram_0_s1_arbitration_holdoff_internal | ~nios_system_clock_5_out_requests_sdram_0_s1) ? 0 : last_cycle_nios_system_clock_5_out_granted_slave_sdram_0_s1;
    end


  //nios_system_clock_5_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_5_out_continuerequest = (last_cycle_nios_system_clock_5_out_granted_slave_sdram_0_s1 & nios_system_clock_5_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_5_out_granted_slave_sdram_0_s1 & nios_system_clock_5_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_5_out_granted_slave_sdram_0_s1 & nios_system_clock_5_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_5_out_granted_slave_sdram_0_s1 & nios_system_clock_5_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_5_out_granted_slave_sdram_0_s1 & nios_system_clock_5_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_5_out_granted_slave_sdram_0_s1 & nios_system_clock_5_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_5_out_granted_slave_sdram_0_s1 & nios_system_clock_5_out_requests_sdram_0_s1);

  //nios_system_clock_6/out sdram_0/s1 arbiterlock, which is an e_assign
  assign nios_system_clock_6_out_arbiterlock = sdram_0_s1_slavearbiterlockenable & nios_system_clock_6_out_continuerequest;

  //nios_system_clock_6/out sdram_0/s1 arbiterlock2, which is an e_assign
  assign nios_system_clock_6_out_arbiterlock2 = sdram_0_s1_slavearbiterlockenable2 & nios_system_clock_6_out_continuerequest;

  //nios_system_clock_6/out granted sdram_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_6_out_granted_slave_sdram_0_s1 <= 0;
      else 
        last_cycle_nios_system_clock_6_out_granted_slave_sdram_0_s1 <= nios_system_clock_6_out_saved_grant_sdram_0_s1 ? 1 : (sdram_0_s1_arbitration_holdoff_internal | ~nios_system_clock_6_out_requests_sdram_0_s1) ? 0 : last_cycle_nios_system_clock_6_out_granted_slave_sdram_0_s1;
    end


  //nios_system_clock_6_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_6_out_continuerequest = (last_cycle_nios_system_clock_6_out_granted_slave_sdram_0_s1 & nios_system_clock_6_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_6_out_granted_slave_sdram_0_s1 & nios_system_clock_6_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_6_out_granted_slave_sdram_0_s1 & nios_system_clock_6_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_6_out_granted_slave_sdram_0_s1 & nios_system_clock_6_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_6_out_granted_slave_sdram_0_s1 & nios_system_clock_6_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_6_out_granted_slave_sdram_0_s1 & nios_system_clock_6_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_6_out_granted_slave_sdram_0_s1 & nios_system_clock_6_out_requests_sdram_0_s1);

  //nios_system_clock_7/out sdram_0/s1 arbiterlock, which is an e_assign
  assign nios_system_clock_7_out_arbiterlock = sdram_0_s1_slavearbiterlockenable & nios_system_clock_7_out_continuerequest;

  //nios_system_clock_7/out sdram_0/s1 arbiterlock2, which is an e_assign
  assign nios_system_clock_7_out_arbiterlock2 = sdram_0_s1_slavearbiterlockenable2 & nios_system_clock_7_out_continuerequest;

  //nios_system_clock_7/out granted sdram_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_7_out_granted_slave_sdram_0_s1 <= 0;
      else 
        last_cycle_nios_system_clock_7_out_granted_slave_sdram_0_s1 <= nios_system_clock_7_out_saved_grant_sdram_0_s1 ? 1 : (sdram_0_s1_arbitration_holdoff_internal | ~nios_system_clock_7_out_requests_sdram_0_s1) ? 0 : last_cycle_nios_system_clock_7_out_granted_slave_sdram_0_s1;
    end


  //nios_system_clock_7_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_7_out_continuerequest = (last_cycle_nios_system_clock_7_out_granted_slave_sdram_0_s1 & nios_system_clock_7_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_7_out_granted_slave_sdram_0_s1 & nios_system_clock_7_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_7_out_granted_slave_sdram_0_s1 & nios_system_clock_7_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_7_out_granted_slave_sdram_0_s1 & nios_system_clock_7_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_7_out_granted_slave_sdram_0_s1 & nios_system_clock_7_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_7_out_granted_slave_sdram_0_s1 & nios_system_clock_7_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_7_out_granted_slave_sdram_0_s1 & nios_system_clock_7_out_requests_sdram_0_s1);

  assign nios_system_clock_0_out_qualified_request_sdram_0_s1 = nios_system_clock_0_out_requests_sdram_0_s1 & ~((nios_system_clock_0_out_read & ((|nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register))) | nios_system_clock_1_out_arbiterlock | nios_system_clock_2_out_arbiterlock | nios_system_clock_3_out_arbiterlock | nios_system_clock_4_out_arbiterlock | nios_system_clock_5_out_arbiterlock | nios_system_clock_6_out_arbiterlock | nios_system_clock_7_out_arbiterlock);
  //unique name for sdram_0_s1_move_on_to_next_transaction, which is an e_assign
  assign sdram_0_s1_move_on_to_next_transaction = sdram_0_s1_readdatavalid_from_sa;

  //rdv_fifo_for_nios_system_clock_0_out_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios_system_clock_0_out_to_sdram_0_s1_module rdv_fifo_for_nios_system_clock_0_out_to_sdram_0_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (nios_system_clock_0_out_granted_sdram_0_s1),
      .data_out             (nios_system_clock_0_out_rdv_fifo_output_from_sdram_0_s1),
      .empty                (),
      .fifo_contains_ones_n (nios_system_clock_0_out_rdv_fifo_empty_sdram_0_s1),
      .full                 (),
      .read                 (sdram_0_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_0_s1_waits_for_read)
    );

  assign nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register = ~nios_system_clock_0_out_rdv_fifo_empty_sdram_0_s1;
  //local readdatavalid nios_system_clock_0_out_read_data_valid_sdram_0_s1, which is an e_mux
  assign nios_system_clock_0_out_read_data_valid_sdram_0_s1 = (sdram_0_s1_readdatavalid_from_sa & nios_system_clock_0_out_rdv_fifo_output_from_sdram_0_s1) & ~ nios_system_clock_0_out_rdv_fifo_empty_sdram_0_s1;

  //sdram_0_s1_writedata mux, which is an e_mux
  assign sdram_0_s1_writedata = (nios_system_clock_0_out_granted_sdram_0_s1)? nios_system_clock_0_out_writedata :
    (nios_system_clock_1_out_granted_sdram_0_s1)? nios_system_clock_1_out_writedata :
    (nios_system_clock_2_out_granted_sdram_0_s1)? nios_system_clock_2_out_writedata :
    (nios_system_clock_3_out_granted_sdram_0_s1)? nios_system_clock_3_out_writedata :
    (nios_system_clock_4_out_granted_sdram_0_s1)? nios_system_clock_4_out_writedata :
    (nios_system_clock_5_out_granted_sdram_0_s1)? nios_system_clock_5_out_writedata :
    (nios_system_clock_6_out_granted_sdram_0_s1)? nios_system_clock_6_out_writedata :
    nios_system_clock_7_out_writedata;

  assign nios_system_clock_1_out_requests_sdram_0_s1 = (1) & (nios_system_clock_1_out_read | nios_system_clock_1_out_write);
  //nios_system_clock_0/out granted sdram_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_nios_system_clock_0_out_granted_slave_sdram_0_s1 <= 0;
      else 
        last_cycle_nios_system_clock_0_out_granted_slave_sdram_0_s1 <= nios_system_clock_0_out_saved_grant_sdram_0_s1 ? 1 : (sdram_0_s1_arbitration_holdoff_internal | ~nios_system_clock_0_out_requests_sdram_0_s1) ? 0 : last_cycle_nios_system_clock_0_out_granted_slave_sdram_0_s1;
    end


  //nios_system_clock_0_out_continuerequest continued request, which is an e_mux
  assign nios_system_clock_0_out_continuerequest = (last_cycle_nios_system_clock_0_out_granted_slave_sdram_0_s1 & nios_system_clock_0_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_0_out_granted_slave_sdram_0_s1 & nios_system_clock_0_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_0_out_granted_slave_sdram_0_s1 & nios_system_clock_0_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_0_out_granted_slave_sdram_0_s1 & nios_system_clock_0_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_0_out_granted_slave_sdram_0_s1 & nios_system_clock_0_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_0_out_granted_slave_sdram_0_s1 & nios_system_clock_0_out_requests_sdram_0_s1) |
    (last_cycle_nios_system_clock_0_out_granted_slave_sdram_0_s1 & nios_system_clock_0_out_requests_sdram_0_s1);

  assign nios_system_clock_1_out_qualified_request_sdram_0_s1 = nios_system_clock_1_out_requests_sdram_0_s1 & ~((nios_system_clock_1_out_read & ((|nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register))) | nios_system_clock_0_out_arbiterlock | nios_system_clock_2_out_arbiterlock | nios_system_clock_3_out_arbiterlock | nios_system_clock_4_out_arbiterlock | nios_system_clock_5_out_arbiterlock | nios_system_clock_6_out_arbiterlock | nios_system_clock_7_out_arbiterlock);
  //rdv_fifo_for_nios_system_clock_1_out_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios_system_clock_1_out_to_sdram_0_s1_module rdv_fifo_for_nios_system_clock_1_out_to_sdram_0_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (nios_system_clock_1_out_granted_sdram_0_s1),
      .data_out             (nios_system_clock_1_out_rdv_fifo_output_from_sdram_0_s1),
      .empty                (),
      .fifo_contains_ones_n (nios_system_clock_1_out_rdv_fifo_empty_sdram_0_s1),
      .full                 (),
      .read                 (sdram_0_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_0_s1_waits_for_read)
    );

  assign nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register = ~nios_system_clock_1_out_rdv_fifo_empty_sdram_0_s1;
  //local readdatavalid nios_system_clock_1_out_read_data_valid_sdram_0_s1, which is an e_mux
  assign nios_system_clock_1_out_read_data_valid_sdram_0_s1 = (sdram_0_s1_readdatavalid_from_sa & nios_system_clock_1_out_rdv_fifo_output_from_sdram_0_s1) & ~ nios_system_clock_1_out_rdv_fifo_empty_sdram_0_s1;

  assign nios_system_clock_2_out_requests_sdram_0_s1 = (1) & (nios_system_clock_2_out_read | nios_system_clock_2_out_write);
  assign nios_system_clock_2_out_qualified_request_sdram_0_s1 = nios_system_clock_2_out_requests_sdram_0_s1 & ~((nios_system_clock_2_out_read & ((|nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register))) | nios_system_clock_0_out_arbiterlock | nios_system_clock_1_out_arbiterlock | nios_system_clock_3_out_arbiterlock | nios_system_clock_4_out_arbiterlock | nios_system_clock_5_out_arbiterlock | nios_system_clock_6_out_arbiterlock | nios_system_clock_7_out_arbiterlock);
  //rdv_fifo_for_nios_system_clock_2_out_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios_system_clock_2_out_to_sdram_0_s1_module rdv_fifo_for_nios_system_clock_2_out_to_sdram_0_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (nios_system_clock_2_out_granted_sdram_0_s1),
      .data_out             (nios_system_clock_2_out_rdv_fifo_output_from_sdram_0_s1),
      .empty                (),
      .fifo_contains_ones_n (nios_system_clock_2_out_rdv_fifo_empty_sdram_0_s1),
      .full                 (),
      .read                 (sdram_0_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_0_s1_waits_for_read)
    );

  assign nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register = ~nios_system_clock_2_out_rdv_fifo_empty_sdram_0_s1;
  //local readdatavalid nios_system_clock_2_out_read_data_valid_sdram_0_s1, which is an e_mux
  assign nios_system_clock_2_out_read_data_valid_sdram_0_s1 = (sdram_0_s1_readdatavalid_from_sa & nios_system_clock_2_out_rdv_fifo_output_from_sdram_0_s1) & ~ nios_system_clock_2_out_rdv_fifo_empty_sdram_0_s1;

  assign nios_system_clock_3_out_requests_sdram_0_s1 = (1) & (nios_system_clock_3_out_read | nios_system_clock_3_out_write);
  assign nios_system_clock_3_out_qualified_request_sdram_0_s1 = nios_system_clock_3_out_requests_sdram_0_s1 & ~((nios_system_clock_3_out_read & ((|nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register))) | nios_system_clock_0_out_arbiterlock | nios_system_clock_1_out_arbiterlock | nios_system_clock_2_out_arbiterlock | nios_system_clock_4_out_arbiterlock | nios_system_clock_5_out_arbiterlock | nios_system_clock_6_out_arbiterlock | nios_system_clock_7_out_arbiterlock);
  //rdv_fifo_for_nios_system_clock_3_out_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios_system_clock_3_out_to_sdram_0_s1_module rdv_fifo_for_nios_system_clock_3_out_to_sdram_0_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (nios_system_clock_3_out_granted_sdram_0_s1),
      .data_out             (nios_system_clock_3_out_rdv_fifo_output_from_sdram_0_s1),
      .empty                (),
      .fifo_contains_ones_n (nios_system_clock_3_out_rdv_fifo_empty_sdram_0_s1),
      .full                 (),
      .read                 (sdram_0_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_0_s1_waits_for_read)
    );

  assign nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register = ~nios_system_clock_3_out_rdv_fifo_empty_sdram_0_s1;
  //local readdatavalid nios_system_clock_3_out_read_data_valid_sdram_0_s1, which is an e_mux
  assign nios_system_clock_3_out_read_data_valid_sdram_0_s1 = (sdram_0_s1_readdatavalid_from_sa & nios_system_clock_3_out_rdv_fifo_output_from_sdram_0_s1) & ~ nios_system_clock_3_out_rdv_fifo_empty_sdram_0_s1;

  assign nios_system_clock_4_out_requests_sdram_0_s1 = (1) & (nios_system_clock_4_out_read | nios_system_clock_4_out_write);
  assign nios_system_clock_4_out_qualified_request_sdram_0_s1 = nios_system_clock_4_out_requests_sdram_0_s1 & ~((nios_system_clock_4_out_read & ((|nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register))) | nios_system_clock_0_out_arbiterlock | nios_system_clock_1_out_arbiterlock | nios_system_clock_2_out_arbiterlock | nios_system_clock_3_out_arbiterlock | nios_system_clock_5_out_arbiterlock | nios_system_clock_6_out_arbiterlock | nios_system_clock_7_out_arbiterlock);
  //rdv_fifo_for_nios_system_clock_4_out_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios_system_clock_4_out_to_sdram_0_s1_module rdv_fifo_for_nios_system_clock_4_out_to_sdram_0_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (nios_system_clock_4_out_granted_sdram_0_s1),
      .data_out             (nios_system_clock_4_out_rdv_fifo_output_from_sdram_0_s1),
      .empty                (),
      .fifo_contains_ones_n (nios_system_clock_4_out_rdv_fifo_empty_sdram_0_s1),
      .full                 (),
      .read                 (sdram_0_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_0_s1_waits_for_read)
    );

  assign nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register = ~nios_system_clock_4_out_rdv_fifo_empty_sdram_0_s1;
  //local readdatavalid nios_system_clock_4_out_read_data_valid_sdram_0_s1, which is an e_mux
  assign nios_system_clock_4_out_read_data_valid_sdram_0_s1 = (sdram_0_s1_readdatavalid_from_sa & nios_system_clock_4_out_rdv_fifo_output_from_sdram_0_s1) & ~ nios_system_clock_4_out_rdv_fifo_empty_sdram_0_s1;

  assign nios_system_clock_5_out_requests_sdram_0_s1 = (1) & (nios_system_clock_5_out_read | nios_system_clock_5_out_write);
  assign nios_system_clock_5_out_qualified_request_sdram_0_s1 = nios_system_clock_5_out_requests_sdram_0_s1 & ~((nios_system_clock_5_out_read & ((|nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register))) | nios_system_clock_0_out_arbiterlock | nios_system_clock_1_out_arbiterlock | nios_system_clock_2_out_arbiterlock | nios_system_clock_3_out_arbiterlock | nios_system_clock_4_out_arbiterlock | nios_system_clock_6_out_arbiterlock | nios_system_clock_7_out_arbiterlock);
  //rdv_fifo_for_nios_system_clock_5_out_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios_system_clock_5_out_to_sdram_0_s1_module rdv_fifo_for_nios_system_clock_5_out_to_sdram_0_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (nios_system_clock_5_out_granted_sdram_0_s1),
      .data_out             (nios_system_clock_5_out_rdv_fifo_output_from_sdram_0_s1),
      .empty                (),
      .fifo_contains_ones_n (nios_system_clock_5_out_rdv_fifo_empty_sdram_0_s1),
      .full                 (),
      .read                 (sdram_0_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_0_s1_waits_for_read)
    );

  assign nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register = ~nios_system_clock_5_out_rdv_fifo_empty_sdram_0_s1;
  //local readdatavalid nios_system_clock_5_out_read_data_valid_sdram_0_s1, which is an e_mux
  assign nios_system_clock_5_out_read_data_valid_sdram_0_s1 = (sdram_0_s1_readdatavalid_from_sa & nios_system_clock_5_out_rdv_fifo_output_from_sdram_0_s1) & ~ nios_system_clock_5_out_rdv_fifo_empty_sdram_0_s1;

  assign nios_system_clock_6_out_requests_sdram_0_s1 = (1) & (nios_system_clock_6_out_read | nios_system_clock_6_out_write);
  assign nios_system_clock_6_out_qualified_request_sdram_0_s1 = nios_system_clock_6_out_requests_sdram_0_s1 & ~((nios_system_clock_6_out_read & ((|nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register))) | nios_system_clock_0_out_arbiterlock | nios_system_clock_1_out_arbiterlock | nios_system_clock_2_out_arbiterlock | nios_system_clock_3_out_arbiterlock | nios_system_clock_4_out_arbiterlock | nios_system_clock_5_out_arbiterlock | nios_system_clock_7_out_arbiterlock);
  //rdv_fifo_for_nios_system_clock_6_out_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios_system_clock_6_out_to_sdram_0_s1_module rdv_fifo_for_nios_system_clock_6_out_to_sdram_0_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (nios_system_clock_6_out_granted_sdram_0_s1),
      .data_out             (nios_system_clock_6_out_rdv_fifo_output_from_sdram_0_s1),
      .empty                (),
      .fifo_contains_ones_n (nios_system_clock_6_out_rdv_fifo_empty_sdram_0_s1),
      .full                 (),
      .read                 (sdram_0_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_0_s1_waits_for_read)
    );

  assign nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register = ~nios_system_clock_6_out_rdv_fifo_empty_sdram_0_s1;
  //local readdatavalid nios_system_clock_6_out_read_data_valid_sdram_0_s1, which is an e_mux
  assign nios_system_clock_6_out_read_data_valid_sdram_0_s1 = (sdram_0_s1_readdatavalid_from_sa & nios_system_clock_6_out_rdv_fifo_output_from_sdram_0_s1) & ~ nios_system_clock_6_out_rdv_fifo_empty_sdram_0_s1;

  assign nios_system_clock_7_out_requests_sdram_0_s1 = (1) & (nios_system_clock_7_out_read | nios_system_clock_7_out_write);
  assign nios_system_clock_7_out_qualified_request_sdram_0_s1 = nios_system_clock_7_out_requests_sdram_0_s1 & ~((nios_system_clock_7_out_read & ((|nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register))) | nios_system_clock_0_out_arbiterlock | nios_system_clock_1_out_arbiterlock | nios_system_clock_2_out_arbiterlock | nios_system_clock_3_out_arbiterlock | nios_system_clock_4_out_arbiterlock | nios_system_clock_5_out_arbiterlock | nios_system_clock_6_out_arbiterlock);
  //rdv_fifo_for_nios_system_clock_7_out_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_nios_system_clock_7_out_to_sdram_0_s1_module rdv_fifo_for_nios_system_clock_7_out_to_sdram_0_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (nios_system_clock_7_out_granted_sdram_0_s1),
      .data_out             (nios_system_clock_7_out_rdv_fifo_output_from_sdram_0_s1),
      .empty                (),
      .fifo_contains_ones_n (nios_system_clock_7_out_rdv_fifo_empty_sdram_0_s1),
      .full                 (),
      .read                 (sdram_0_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_0_s1_waits_for_read)
    );

  assign nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register = ~nios_system_clock_7_out_rdv_fifo_empty_sdram_0_s1;
  //local readdatavalid nios_system_clock_7_out_read_data_valid_sdram_0_s1, which is an e_mux
  assign nios_system_clock_7_out_read_data_valid_sdram_0_s1 = (sdram_0_s1_readdatavalid_from_sa & nios_system_clock_7_out_rdv_fifo_output_from_sdram_0_s1) & ~ nios_system_clock_7_out_rdv_fifo_empty_sdram_0_s1;

  //allow new arb cycle for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_allow_new_arb_cycle = ~nios_system_clock_0_out_arbiterlock & ~nios_system_clock_1_out_arbiterlock & ~nios_system_clock_2_out_arbiterlock & ~nios_system_clock_3_out_arbiterlock & ~nios_system_clock_4_out_arbiterlock & ~nios_system_clock_5_out_arbiterlock & ~nios_system_clock_6_out_arbiterlock & ~nios_system_clock_7_out_arbiterlock;

  //nios_system_clock_7/out assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_master_qreq_vector[0] = nios_system_clock_7_out_qualified_request_sdram_0_s1;

  //nios_system_clock_7/out grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_7_out_granted_sdram_0_s1 = sdram_0_s1_grant_vector[0];

  //nios_system_clock_7/out saved-grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_7_out_saved_grant_sdram_0_s1 = sdram_0_s1_arb_winner[0] && nios_system_clock_7_out_requests_sdram_0_s1;

  //nios_system_clock_6/out assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_master_qreq_vector[1] = nios_system_clock_6_out_qualified_request_sdram_0_s1;

  //nios_system_clock_6/out grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_6_out_granted_sdram_0_s1 = sdram_0_s1_grant_vector[1];

  //nios_system_clock_6/out saved-grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_6_out_saved_grant_sdram_0_s1 = sdram_0_s1_arb_winner[1] && nios_system_clock_6_out_requests_sdram_0_s1;

  //nios_system_clock_5/out assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_master_qreq_vector[2] = nios_system_clock_5_out_qualified_request_sdram_0_s1;

  //nios_system_clock_5/out grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_5_out_granted_sdram_0_s1 = sdram_0_s1_grant_vector[2];

  //nios_system_clock_5/out saved-grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_5_out_saved_grant_sdram_0_s1 = sdram_0_s1_arb_winner[2] && nios_system_clock_5_out_requests_sdram_0_s1;

  //nios_system_clock_4/out assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_master_qreq_vector[3] = nios_system_clock_4_out_qualified_request_sdram_0_s1;

  //nios_system_clock_4/out grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_4_out_granted_sdram_0_s1 = sdram_0_s1_grant_vector[3];

  //nios_system_clock_4/out saved-grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_4_out_saved_grant_sdram_0_s1 = sdram_0_s1_arb_winner[3] && nios_system_clock_4_out_requests_sdram_0_s1;

  //nios_system_clock_3/out assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_master_qreq_vector[4] = nios_system_clock_3_out_qualified_request_sdram_0_s1;

  //nios_system_clock_3/out grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_3_out_granted_sdram_0_s1 = sdram_0_s1_grant_vector[4];

  //nios_system_clock_3/out saved-grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_3_out_saved_grant_sdram_0_s1 = sdram_0_s1_arb_winner[4] && nios_system_clock_3_out_requests_sdram_0_s1;

  //nios_system_clock_2/out assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_master_qreq_vector[5] = nios_system_clock_2_out_qualified_request_sdram_0_s1;

  //nios_system_clock_2/out grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_2_out_granted_sdram_0_s1 = sdram_0_s1_grant_vector[5];

  //nios_system_clock_2/out saved-grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_2_out_saved_grant_sdram_0_s1 = sdram_0_s1_arb_winner[5] && nios_system_clock_2_out_requests_sdram_0_s1;

  //nios_system_clock_1/out assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_master_qreq_vector[6] = nios_system_clock_1_out_qualified_request_sdram_0_s1;

  //nios_system_clock_1/out grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_1_out_granted_sdram_0_s1 = sdram_0_s1_grant_vector[6];

  //nios_system_clock_1/out saved-grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_1_out_saved_grant_sdram_0_s1 = sdram_0_s1_arb_winner[6] && nios_system_clock_1_out_requests_sdram_0_s1;

  //nios_system_clock_0/out assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_master_qreq_vector[7] = nios_system_clock_0_out_qualified_request_sdram_0_s1;

  //nios_system_clock_0/out grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_0_out_granted_sdram_0_s1 = sdram_0_s1_grant_vector[7];

  //nios_system_clock_0/out saved-grant sdram_0/s1, which is an e_assign
  assign nios_system_clock_0_out_saved_grant_sdram_0_s1 = sdram_0_s1_arb_winner[7] && nios_system_clock_0_out_requests_sdram_0_s1;

  //sdram_0/s1 chosen-master double-vector, which is an e_assign
  assign sdram_0_s1_chosen_master_double_vector = {sdram_0_s1_master_qreq_vector, sdram_0_s1_master_qreq_vector} & ({~sdram_0_s1_master_qreq_vector, ~sdram_0_s1_master_qreq_vector} + sdram_0_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign sdram_0_s1_arb_winner = (sdram_0_s1_allow_new_arb_cycle & | sdram_0_s1_grant_vector) ? sdram_0_s1_grant_vector : sdram_0_s1_saved_chosen_master_vector;

  //saved sdram_0_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_0_s1_saved_chosen_master_vector <= 0;
      else if (sdram_0_s1_allow_new_arb_cycle)
          sdram_0_s1_saved_chosen_master_vector <= |sdram_0_s1_grant_vector ? sdram_0_s1_grant_vector : sdram_0_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign sdram_0_s1_grant_vector = {(sdram_0_s1_chosen_master_double_vector[7] | sdram_0_s1_chosen_master_double_vector[15]),
    (sdram_0_s1_chosen_master_double_vector[6] | sdram_0_s1_chosen_master_double_vector[14]),
    (sdram_0_s1_chosen_master_double_vector[5] | sdram_0_s1_chosen_master_double_vector[13]),
    (sdram_0_s1_chosen_master_double_vector[4] | sdram_0_s1_chosen_master_double_vector[12]),
    (sdram_0_s1_chosen_master_double_vector[3] | sdram_0_s1_chosen_master_double_vector[11]),
    (sdram_0_s1_chosen_master_double_vector[2] | sdram_0_s1_chosen_master_double_vector[10]),
    (sdram_0_s1_chosen_master_double_vector[1] | sdram_0_s1_chosen_master_double_vector[9]),
    (sdram_0_s1_chosen_master_double_vector[0] | sdram_0_s1_chosen_master_double_vector[8])};

  //sdram_0/s1 chosen master rotated left, which is an e_assign
  assign sdram_0_s1_chosen_master_rot_left = (sdram_0_s1_arb_winner << 1) ? (sdram_0_s1_arb_winner << 1) : 1;

  //sdram_0/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_0_s1_arb_addend <= 1;
      else if (|sdram_0_s1_grant_vector)
          sdram_0_s1_arb_addend <= sdram_0_s1_end_xfer? sdram_0_s1_chosen_master_rot_left : sdram_0_s1_grant_vector;
    end


  //sdram_0_s1_reset_n assignment, which is an e_assign
  assign sdram_0_s1_reset_n = reset_n;

  assign sdram_0_s1_chipselect = nios_system_clock_0_out_granted_sdram_0_s1 | nios_system_clock_1_out_granted_sdram_0_s1 | nios_system_clock_2_out_granted_sdram_0_s1 | nios_system_clock_3_out_granted_sdram_0_s1 | nios_system_clock_4_out_granted_sdram_0_s1 | nios_system_clock_5_out_granted_sdram_0_s1 | nios_system_clock_6_out_granted_sdram_0_s1 | nios_system_clock_7_out_granted_sdram_0_s1;
  //sdram_0_s1_firsttransfer first transaction, which is an e_assign
  assign sdram_0_s1_firsttransfer = sdram_0_s1_begins_xfer ? sdram_0_s1_unreg_firsttransfer : sdram_0_s1_reg_firsttransfer;

  //sdram_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign sdram_0_s1_unreg_firsttransfer = ~(sdram_0_s1_slavearbiterlockenable & sdram_0_s1_any_continuerequest);

  //sdram_0_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_0_s1_reg_firsttransfer <= 1'b1;
      else if (sdram_0_s1_begins_xfer)
          sdram_0_s1_reg_firsttransfer <= sdram_0_s1_unreg_firsttransfer;
    end


  //sdram_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sdram_0_s1_beginbursttransfer_internal = sdram_0_s1_begins_xfer;

  //sdram_0_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign sdram_0_s1_arbitration_holdoff_internal = sdram_0_s1_begins_xfer & sdram_0_s1_firsttransfer;

  //~sdram_0_s1_read_n assignment, which is an e_mux
  assign sdram_0_s1_read_n = ~((nios_system_clock_0_out_granted_sdram_0_s1 & nios_system_clock_0_out_read) | (nios_system_clock_1_out_granted_sdram_0_s1 & nios_system_clock_1_out_read) | (nios_system_clock_2_out_granted_sdram_0_s1 & nios_system_clock_2_out_read) | (nios_system_clock_3_out_granted_sdram_0_s1 & nios_system_clock_3_out_read) | (nios_system_clock_4_out_granted_sdram_0_s1 & nios_system_clock_4_out_read) | (nios_system_clock_5_out_granted_sdram_0_s1 & nios_system_clock_5_out_read) | (nios_system_clock_6_out_granted_sdram_0_s1 & nios_system_clock_6_out_read) | (nios_system_clock_7_out_granted_sdram_0_s1 & nios_system_clock_7_out_read));

  //~sdram_0_s1_write_n assignment, which is an e_mux
  assign sdram_0_s1_write_n = ~((nios_system_clock_0_out_granted_sdram_0_s1 & nios_system_clock_0_out_write) | (nios_system_clock_1_out_granted_sdram_0_s1 & nios_system_clock_1_out_write) | (nios_system_clock_2_out_granted_sdram_0_s1 & nios_system_clock_2_out_write) | (nios_system_clock_3_out_granted_sdram_0_s1 & nios_system_clock_3_out_write) | (nios_system_clock_4_out_granted_sdram_0_s1 & nios_system_clock_4_out_write) | (nios_system_clock_5_out_granted_sdram_0_s1 & nios_system_clock_5_out_write) | (nios_system_clock_6_out_granted_sdram_0_s1 & nios_system_clock_6_out_write) | (nios_system_clock_7_out_granted_sdram_0_s1 & nios_system_clock_7_out_write));

  assign shifted_address_to_sdram_0_s1_from_nios_system_clock_0_out = nios_system_clock_0_out_address_to_slave;
  //sdram_0_s1_address mux, which is an e_mux
  assign sdram_0_s1_address = (nios_system_clock_0_out_granted_sdram_0_s1)? (shifted_address_to_sdram_0_s1_from_nios_system_clock_0_out >> 1) :
    (nios_system_clock_1_out_granted_sdram_0_s1)? (shifted_address_to_sdram_0_s1_from_nios_system_clock_1_out >> 1) :
    (nios_system_clock_2_out_granted_sdram_0_s1)? (shifted_address_to_sdram_0_s1_from_nios_system_clock_2_out >> 1) :
    (nios_system_clock_3_out_granted_sdram_0_s1)? (shifted_address_to_sdram_0_s1_from_nios_system_clock_3_out >> 1) :
    (nios_system_clock_4_out_granted_sdram_0_s1)? (shifted_address_to_sdram_0_s1_from_nios_system_clock_4_out >> 1) :
    (nios_system_clock_5_out_granted_sdram_0_s1)? (shifted_address_to_sdram_0_s1_from_nios_system_clock_5_out >> 1) :
    (nios_system_clock_6_out_granted_sdram_0_s1)? (shifted_address_to_sdram_0_s1_from_nios_system_clock_6_out >> 1) :
    (shifted_address_to_sdram_0_s1_from_nios_system_clock_7_out >> 1);

  assign shifted_address_to_sdram_0_s1_from_nios_system_clock_1_out = nios_system_clock_1_out_address_to_slave;
  assign shifted_address_to_sdram_0_s1_from_nios_system_clock_2_out = nios_system_clock_2_out_address_to_slave;
  assign shifted_address_to_sdram_0_s1_from_nios_system_clock_3_out = nios_system_clock_3_out_address_to_slave;
  assign shifted_address_to_sdram_0_s1_from_nios_system_clock_4_out = nios_system_clock_4_out_address_to_slave;
  assign shifted_address_to_sdram_0_s1_from_nios_system_clock_5_out = nios_system_clock_5_out_address_to_slave;
  assign shifted_address_to_sdram_0_s1_from_nios_system_clock_6_out = nios_system_clock_6_out_address_to_slave;
  assign shifted_address_to_sdram_0_s1_from_nios_system_clock_7_out = nios_system_clock_7_out_address_to_slave;
  //d1_sdram_0_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sdram_0_s1_end_xfer <= 1;
      else 
        d1_sdram_0_s1_end_xfer <= sdram_0_s1_end_xfer;
    end


  //sdram_0_s1_waits_for_read in a cycle, which is an e_mux
  assign sdram_0_s1_waits_for_read = sdram_0_s1_in_a_read_cycle & sdram_0_s1_waitrequest_from_sa;

  //sdram_0_s1_in_a_read_cycle assignment, which is an e_assign
  assign sdram_0_s1_in_a_read_cycle = (nios_system_clock_0_out_granted_sdram_0_s1 & nios_system_clock_0_out_read) | (nios_system_clock_1_out_granted_sdram_0_s1 & nios_system_clock_1_out_read) | (nios_system_clock_2_out_granted_sdram_0_s1 & nios_system_clock_2_out_read) | (nios_system_clock_3_out_granted_sdram_0_s1 & nios_system_clock_3_out_read) | (nios_system_clock_4_out_granted_sdram_0_s1 & nios_system_clock_4_out_read) | (nios_system_clock_5_out_granted_sdram_0_s1 & nios_system_clock_5_out_read) | (nios_system_clock_6_out_granted_sdram_0_s1 & nios_system_clock_6_out_read) | (nios_system_clock_7_out_granted_sdram_0_s1 & nios_system_clock_7_out_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sdram_0_s1_in_a_read_cycle;

  //sdram_0_s1_waits_for_write in a cycle, which is an e_mux
  assign sdram_0_s1_waits_for_write = sdram_0_s1_in_a_write_cycle & sdram_0_s1_waitrequest_from_sa;

  //sdram_0_s1_in_a_write_cycle assignment, which is an e_assign
  assign sdram_0_s1_in_a_write_cycle = (nios_system_clock_0_out_granted_sdram_0_s1 & nios_system_clock_0_out_write) | (nios_system_clock_1_out_granted_sdram_0_s1 & nios_system_clock_1_out_write) | (nios_system_clock_2_out_granted_sdram_0_s1 & nios_system_clock_2_out_write) | (nios_system_clock_3_out_granted_sdram_0_s1 & nios_system_clock_3_out_write) | (nios_system_clock_4_out_granted_sdram_0_s1 & nios_system_clock_4_out_write) | (nios_system_clock_5_out_granted_sdram_0_s1 & nios_system_clock_5_out_write) | (nios_system_clock_6_out_granted_sdram_0_s1 & nios_system_clock_6_out_write) | (nios_system_clock_7_out_granted_sdram_0_s1 & nios_system_clock_7_out_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sdram_0_s1_in_a_write_cycle;

  assign wait_for_sdram_0_s1_counter = 0;
  //~sdram_0_s1_byteenable_n byte enable port mux, which is an e_mux
  assign sdram_0_s1_byteenable_n = ~((nios_system_clock_0_out_granted_sdram_0_s1)? nios_system_clock_0_out_byteenable :
    (nios_system_clock_1_out_granted_sdram_0_s1)? nios_system_clock_1_out_byteenable :
    (nios_system_clock_2_out_granted_sdram_0_s1)? nios_system_clock_2_out_byteenable :
    (nios_system_clock_3_out_granted_sdram_0_s1)? nios_system_clock_3_out_byteenable :
    (nios_system_clock_4_out_granted_sdram_0_s1)? nios_system_clock_4_out_byteenable :
    (nios_system_clock_5_out_granted_sdram_0_s1)? nios_system_clock_5_out_byteenable :
    (nios_system_clock_6_out_granted_sdram_0_s1)? nios_system_clock_6_out_byteenable :
    (nios_system_clock_7_out_granted_sdram_0_s1)? nios_system_clock_7_out_byteenable :
    -1);


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sdram_0/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (nios_system_clock_0_out_granted_sdram_0_s1 + nios_system_clock_1_out_granted_sdram_0_s1 + nios_system_clock_2_out_granted_sdram_0_s1 + nios_system_clock_3_out_granted_sdram_0_s1 + nios_system_clock_4_out_granted_sdram_0_s1 + nios_system_clock_5_out_granted_sdram_0_s1 + nios_system_clock_6_out_granted_sdram_0_s1 + nios_system_clock_7_out_granted_sdram_0_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (nios_system_clock_0_out_saved_grant_sdram_0_s1 + nios_system_clock_1_out_saved_grant_sdram_0_s1 + nios_system_clock_2_out_saved_grant_sdram_0_s1 + nios_system_clock_3_out_saved_grant_sdram_0_s1 + nios_system_clock_4_out_saved_grant_sdram_0_s1 + nios_system_clock_5_out_saved_grant_sdram_0_s1 + nios_system_clock_6_out_saved_grant_sdram_0_s1 + nios_system_clock_7_out_saved_grant_sdram_0_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_0_data_master_to_sram_0_avalon_sram_slave_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_1_data_master_to_sram_0_avalon_sram_slave_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_1_instruction_master_to_sram_0_avalon_sram_slave_module (
                                                                                  // inputs:
                                                                                   clear_fifo,
                                                                                   clk,
                                                                                   data_in,
                                                                                   read,
                                                                                   reset_n,
                                                                                   sync_reset,
                                                                                   write,

                                                                                  // outputs:
                                                                                   data_out,
                                                                                   empty,
                                                                                   fifo_contains_ones_n,
                                                                                   full
                                                                                )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_2_data_master_to_sram_0_avalon_sram_slave_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_2_instruction_master_to_sram_0_avalon_sram_slave_module (
                                                                                  // inputs:
                                                                                   clear_fifo,
                                                                                   clk,
                                                                                   data_in,
                                                                                   read,
                                                                                   reset_n,
                                                                                   sync_reset,
                                                                                   write,

                                                                                  // outputs:
                                                                                   data_out,
                                                                                   empty,
                                                                                   fifo_contains_ones_n,
                                                                                   full
                                                                                )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_3_data_master_to_sram_0_avalon_sram_slave_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_3_instruction_master_to_sram_0_avalon_sram_slave_module (
                                                                                  // inputs:
                                                                                   clear_fifo,
                                                                                   clk,
                                                                                   data_in,
                                                                                   read,
                                                                                   reset_n,
                                                                                   sync_reset,
                                                                                   write,

                                                                                  // outputs:
                                                                                   data_out,
                                                                                   empty,
                                                                                   fifo_contains_ones_n,
                                                                                   full
                                                                                )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_video_pixel_buffer_dma_0_avalon_pixel_dma_master_to_sram_0_avalon_sram_slave_module (
                                                                                                          // inputs:
                                                                                                           clear_fifo,
                                                                                                           clk,
                                                                                                           data_in,
                                                                                                           read,
                                                                                                           reset_n,
                                                                                                           sync_reset,
                                                                                                           write,

                                                                                                          // outputs:
                                                                                                           data_out,
                                                                                                           empty,
                                                                                                           fifo_contains_ones_n,
                                                                                                           full
                                                                                                        )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  wire             full_2;
  reg     [  2: 0] how_many_ones;
  wire    [  2: 0] one_count_minus_one;
  wire    [  2: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  reg              stage_0;
  reg              stage_1;
  wire    [  2: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_1;
  assign empty = !full_0;
  assign full_2 = 0;
  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    0;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sram_0_avalon_sram_slave_arbitrator (
                                             // inputs:
                                              clk,
                                              cpu_0_data_master_address_to_slave,
                                              cpu_0_data_master_byteenable,
                                              cpu_0_data_master_dbs_address,
                                              cpu_0_data_master_dbs_write_16,
                                              cpu_0_data_master_latency_counter,
                                              cpu_0_data_master_read,
                                              cpu_0_data_master_write,
                                              cpu_1_data_master_address_to_slave,
                                              cpu_1_data_master_byteenable,
                                              cpu_1_data_master_dbs_address,
                                              cpu_1_data_master_dbs_write_16,
                                              cpu_1_data_master_latency_counter,
                                              cpu_1_data_master_read,
                                              cpu_1_data_master_write,
                                              cpu_1_instruction_master_address_to_slave,
                                              cpu_1_instruction_master_dbs_address,
                                              cpu_1_instruction_master_latency_counter,
                                              cpu_1_instruction_master_read,
                                              cpu_2_data_master_address_to_slave,
                                              cpu_2_data_master_byteenable,
                                              cpu_2_data_master_dbs_address,
                                              cpu_2_data_master_dbs_write_16,
                                              cpu_2_data_master_latency_counter,
                                              cpu_2_data_master_read,
                                              cpu_2_data_master_write,
                                              cpu_2_instruction_master_address_to_slave,
                                              cpu_2_instruction_master_dbs_address,
                                              cpu_2_instruction_master_latency_counter,
                                              cpu_2_instruction_master_read,
                                              cpu_3_data_master_address_to_slave,
                                              cpu_3_data_master_byteenable,
                                              cpu_3_data_master_dbs_address,
                                              cpu_3_data_master_dbs_write_16,
                                              cpu_3_data_master_latency_counter,
                                              cpu_3_data_master_read,
                                              cpu_3_data_master_write,
                                              cpu_3_instruction_master_address_to_slave,
                                              cpu_3_instruction_master_dbs_address,
                                              cpu_3_instruction_master_latency_counter,
                                              cpu_3_instruction_master_read,
                                              reset_n,
                                              sram_0_avalon_sram_slave_readdata,
                                              sram_0_avalon_sram_slave_readdatavalid,
                                              video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave,
                                              video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock,
                                              video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address,
                                              video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter,
                                              video_pixel_buffer_dma_0_avalon_pixel_dma_master_read,

                                             // outputs:
                                              cpu_0_data_master_byteenable_sram_0_avalon_sram_slave,
                                              cpu_0_data_master_granted_sram_0_avalon_sram_slave,
                                              cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave,
                                              cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave,
                                              cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                              cpu_0_data_master_requests_sram_0_avalon_sram_slave,
                                              cpu_1_data_master_byteenable_sram_0_avalon_sram_slave,
                                              cpu_1_data_master_granted_sram_0_avalon_sram_slave,
                                              cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave,
                                              cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave,
                                              cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                              cpu_1_data_master_requests_sram_0_avalon_sram_slave,
                                              cpu_1_instruction_master_granted_sram_0_avalon_sram_slave,
                                              cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave,
                                              cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave,
                                              cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                              cpu_1_instruction_master_requests_sram_0_avalon_sram_slave,
                                              cpu_2_data_master_byteenable_sram_0_avalon_sram_slave,
                                              cpu_2_data_master_granted_sram_0_avalon_sram_slave,
                                              cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave,
                                              cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave,
                                              cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                              cpu_2_data_master_requests_sram_0_avalon_sram_slave,
                                              cpu_2_instruction_master_granted_sram_0_avalon_sram_slave,
                                              cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave,
                                              cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave,
                                              cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                              cpu_2_instruction_master_requests_sram_0_avalon_sram_slave,
                                              cpu_3_data_master_byteenable_sram_0_avalon_sram_slave,
                                              cpu_3_data_master_granted_sram_0_avalon_sram_slave,
                                              cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave,
                                              cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave,
                                              cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                              cpu_3_data_master_requests_sram_0_avalon_sram_slave,
                                              cpu_3_instruction_master_granted_sram_0_avalon_sram_slave,
                                              cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave,
                                              cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave,
                                              cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                              cpu_3_instruction_master_requests_sram_0_avalon_sram_slave,
                                              d1_sram_0_avalon_sram_slave_end_xfer,
                                              sram_0_avalon_sram_slave_address,
                                              sram_0_avalon_sram_slave_byteenable,
                                              sram_0_avalon_sram_slave_read,
                                              sram_0_avalon_sram_slave_readdata_from_sa,
                                              sram_0_avalon_sram_slave_reset,
                                              sram_0_avalon_sram_slave_write,
                                              sram_0_avalon_sram_slave_writedata,
                                              video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave,
                                              video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave,
                                              video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave,
                                              video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                              video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave
                                           )
;

  output  [  1: 0] cpu_0_data_master_byteenable_sram_0_avalon_sram_slave;
  output           cpu_0_data_master_granted_sram_0_avalon_sram_slave;
  output           cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave;
  output           cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave;
  output           cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  output           cpu_0_data_master_requests_sram_0_avalon_sram_slave;
  output  [  1: 0] cpu_1_data_master_byteenable_sram_0_avalon_sram_slave;
  output           cpu_1_data_master_granted_sram_0_avalon_sram_slave;
  output           cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave;
  output           cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave;
  output           cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  output           cpu_1_data_master_requests_sram_0_avalon_sram_slave;
  output           cpu_1_instruction_master_granted_sram_0_avalon_sram_slave;
  output           cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  output           cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  output           cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  output           cpu_1_instruction_master_requests_sram_0_avalon_sram_slave;
  output  [  1: 0] cpu_2_data_master_byteenable_sram_0_avalon_sram_slave;
  output           cpu_2_data_master_granted_sram_0_avalon_sram_slave;
  output           cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave;
  output           cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave;
  output           cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  output           cpu_2_data_master_requests_sram_0_avalon_sram_slave;
  output           cpu_2_instruction_master_granted_sram_0_avalon_sram_slave;
  output           cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  output           cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  output           cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  output           cpu_2_instruction_master_requests_sram_0_avalon_sram_slave;
  output  [  1: 0] cpu_3_data_master_byteenable_sram_0_avalon_sram_slave;
  output           cpu_3_data_master_granted_sram_0_avalon_sram_slave;
  output           cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave;
  output           cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave;
  output           cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  output           cpu_3_data_master_requests_sram_0_avalon_sram_slave;
  output           cpu_3_instruction_master_granted_sram_0_avalon_sram_slave;
  output           cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  output           cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  output           cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  output           cpu_3_instruction_master_requests_sram_0_avalon_sram_slave;
  output           d1_sram_0_avalon_sram_slave_end_xfer;
  output  [ 17: 0] sram_0_avalon_sram_slave_address;
  output  [  1: 0] sram_0_avalon_sram_slave_byteenable;
  output           sram_0_avalon_sram_slave_read;
  output  [ 15: 0] sram_0_avalon_sram_slave_readdata_from_sa;
  output           sram_0_avalon_sram_slave_reset;
  output           sram_0_avalon_sram_slave_write;
  output  [ 15: 0] sram_0_avalon_sram_slave_writedata;
  output           video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave;
  output           video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave;
  output           video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave;
  output           video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  output           video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input   [  1: 0] cpu_0_data_master_dbs_address;
  input   [ 15: 0] cpu_0_data_master_dbs_write_16;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_write;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input   [  3: 0] cpu_1_data_master_byteenable;
  input   [  1: 0] cpu_1_data_master_dbs_address;
  input   [ 15: 0] cpu_1_data_master_dbs_write_16;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_write;
  input   [ 24: 0] cpu_1_instruction_master_address_to_slave;
  input   [  1: 0] cpu_1_instruction_master_dbs_address;
  input            cpu_1_instruction_master_latency_counter;
  input            cpu_1_instruction_master_read;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input   [  3: 0] cpu_2_data_master_byteenable;
  input   [  1: 0] cpu_2_data_master_dbs_address;
  input   [ 15: 0] cpu_2_data_master_dbs_write_16;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_write;
  input   [ 24: 0] cpu_2_instruction_master_address_to_slave;
  input   [  1: 0] cpu_2_instruction_master_dbs_address;
  input            cpu_2_instruction_master_latency_counter;
  input            cpu_2_instruction_master_read;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input   [  3: 0] cpu_3_data_master_byteenable;
  input   [  1: 0] cpu_3_data_master_dbs_address;
  input   [ 15: 0] cpu_3_data_master_dbs_write_16;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_write;
  input   [ 24: 0] cpu_3_instruction_master_address_to_slave;
  input   [  1: 0] cpu_3_instruction_master_dbs_address;
  input            cpu_3_instruction_master_latency_counter;
  input            cpu_3_instruction_master_read;
  input            reset_n;
  input   [ 15: 0] sram_0_avalon_sram_slave_readdata;
  input            sram_0_avalon_sram_slave_readdatavalid;
  input   [ 31: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave;
  input            video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock;
  input   [  1: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address;
  input            video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter;
  input            video_pixel_buffer_dma_0_avalon_pixel_dma_master_read;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire    [  1: 0] cpu_0_data_master_byteenable_sram_0_avalon_sram_slave;
  wire    [  1: 0] cpu_0_data_master_byteenable_sram_0_avalon_sram_slave_segment_0;
  wire    [  1: 0] cpu_0_data_master_byteenable_sram_0_avalon_sram_slave_segment_1;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_0_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  wire             cpu_0_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave;
  wire             cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             cpu_0_data_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_0_data_master_saved_grant_sram_0_avalon_sram_slave;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire    [  1: 0] cpu_1_data_master_byteenable_sram_0_avalon_sram_slave;
  wire    [  1: 0] cpu_1_data_master_byteenable_sram_0_avalon_sram_slave_segment_0;
  wire    [  1: 0] cpu_1_data_master_byteenable_sram_0_avalon_sram_slave_segment_1;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_1_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  wire             cpu_1_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave;
  wire             cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             cpu_1_data_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_1_data_master_saved_grant_sram_0_avalon_sram_slave;
  wire             cpu_1_instruction_master_arbiterlock;
  wire             cpu_1_instruction_master_arbiterlock2;
  wire             cpu_1_instruction_master_continuerequest;
  wire             cpu_1_instruction_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_1_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  wire             cpu_1_instruction_master_rdv_fifo_output_from_sram_0_avalon_sram_slave;
  wire             cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             cpu_1_instruction_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_1_instruction_master_saved_grant_sram_0_avalon_sram_slave;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire    [  1: 0] cpu_2_data_master_byteenable_sram_0_avalon_sram_slave;
  wire    [  1: 0] cpu_2_data_master_byteenable_sram_0_avalon_sram_slave_segment_0;
  wire    [  1: 0] cpu_2_data_master_byteenable_sram_0_avalon_sram_slave_segment_1;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_2_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  wire             cpu_2_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave;
  wire             cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             cpu_2_data_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_2_data_master_saved_grant_sram_0_avalon_sram_slave;
  wire             cpu_2_instruction_master_arbiterlock;
  wire             cpu_2_instruction_master_arbiterlock2;
  wire             cpu_2_instruction_master_continuerequest;
  wire             cpu_2_instruction_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_2_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  wire             cpu_2_instruction_master_rdv_fifo_output_from_sram_0_avalon_sram_slave;
  wire             cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             cpu_2_instruction_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_2_instruction_master_saved_grant_sram_0_avalon_sram_slave;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire    [  1: 0] cpu_3_data_master_byteenable_sram_0_avalon_sram_slave;
  wire    [  1: 0] cpu_3_data_master_byteenable_sram_0_avalon_sram_slave_segment_0;
  wire    [  1: 0] cpu_3_data_master_byteenable_sram_0_avalon_sram_slave_segment_1;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_3_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  wire             cpu_3_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave;
  wire             cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             cpu_3_data_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_3_data_master_saved_grant_sram_0_avalon_sram_slave;
  wire             cpu_3_instruction_master_arbiterlock;
  wire             cpu_3_instruction_master_arbiterlock2;
  wire             cpu_3_instruction_master_continuerequest;
  wire             cpu_3_instruction_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_3_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  wire             cpu_3_instruction_master_rdv_fifo_output_from_sram_0_avalon_sram_slave;
  wire             cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             cpu_3_instruction_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_3_instruction_master_saved_grant_sram_0_avalon_sram_slave;
  reg              d1_reasons_to_wait;
  reg              d1_sram_0_avalon_sram_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sram_0_avalon_sram_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_sram_0_avalon_sram_slave;
  reg              last_cycle_cpu_1_data_master_granted_slave_sram_0_avalon_sram_slave;
  reg              last_cycle_cpu_1_instruction_master_granted_slave_sram_0_avalon_sram_slave;
  reg              last_cycle_cpu_2_data_master_granted_slave_sram_0_avalon_sram_slave;
  reg              last_cycle_cpu_2_instruction_master_granted_slave_sram_0_avalon_sram_slave;
  reg              last_cycle_cpu_3_data_master_granted_slave_sram_0_avalon_sram_slave;
  reg              last_cycle_cpu_3_instruction_master_granted_slave_sram_0_avalon_sram_slave;
  reg              last_cycle_video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_slave_sram_0_avalon_sram_slave;
  wire             saved_chosen_master_btw_video_pixel_buffer_dma_0_avalon_pixel_dma_master_and_sram_0_avalon_sram_slave;
  wire    [ 24: 0] shifted_address_to_sram_0_avalon_sram_slave_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_sram_0_avalon_sram_slave_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_sram_0_avalon_sram_slave_from_cpu_1_instruction_master;
  wire    [ 24: 0] shifted_address_to_sram_0_avalon_sram_slave_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_sram_0_avalon_sram_slave_from_cpu_2_instruction_master;
  wire    [ 24: 0] shifted_address_to_sram_0_avalon_sram_slave_from_cpu_3_data_master;
  wire    [ 24: 0] shifted_address_to_sram_0_avalon_sram_slave_from_cpu_3_instruction_master;
  wire    [ 31: 0] shifted_address_to_sram_0_avalon_sram_slave_from_video_pixel_buffer_dma_0_avalon_pixel_dma_master;
  wire    [ 17: 0] sram_0_avalon_sram_slave_address;
  wire             sram_0_avalon_sram_slave_allgrants;
  wire             sram_0_avalon_sram_slave_allow_new_arb_cycle;
  wire             sram_0_avalon_sram_slave_any_bursting_master_saved_grant;
  wire             sram_0_avalon_sram_slave_any_continuerequest;
  reg     [  7: 0] sram_0_avalon_sram_slave_arb_addend;
  wire             sram_0_avalon_sram_slave_arb_counter_enable;
  reg     [  2: 0] sram_0_avalon_sram_slave_arb_share_counter;
  wire    [  2: 0] sram_0_avalon_sram_slave_arb_share_counter_next_value;
  wire    [  2: 0] sram_0_avalon_sram_slave_arb_share_set_values;
  wire    [  7: 0] sram_0_avalon_sram_slave_arb_winner;
  wire             sram_0_avalon_sram_slave_arbitration_holdoff_internal;
  wire             sram_0_avalon_sram_slave_beginbursttransfer_internal;
  wire             sram_0_avalon_sram_slave_begins_xfer;
  wire    [  1: 0] sram_0_avalon_sram_slave_byteenable;
  wire    [ 15: 0] sram_0_avalon_sram_slave_chosen_master_double_vector;
  wire    [  7: 0] sram_0_avalon_sram_slave_chosen_master_rot_left;
  wire             sram_0_avalon_sram_slave_end_xfer;
  wire             sram_0_avalon_sram_slave_firsttransfer;
  wire    [  7: 0] sram_0_avalon_sram_slave_grant_vector;
  wire             sram_0_avalon_sram_slave_in_a_read_cycle;
  wire             sram_0_avalon_sram_slave_in_a_write_cycle;
  wire    [  7: 0] sram_0_avalon_sram_slave_master_qreq_vector;
  wire             sram_0_avalon_sram_slave_move_on_to_next_transaction;
  wire             sram_0_avalon_sram_slave_non_bursting_master_requests;
  wire             sram_0_avalon_sram_slave_read;
  wire    [ 15: 0] sram_0_avalon_sram_slave_readdata_from_sa;
  wire             sram_0_avalon_sram_slave_readdatavalid_from_sa;
  reg              sram_0_avalon_sram_slave_reg_firsttransfer;
  wire             sram_0_avalon_sram_slave_reset;
  reg     [  7: 0] sram_0_avalon_sram_slave_saved_chosen_master_vector;
  reg              sram_0_avalon_sram_slave_slavearbiterlockenable;
  wire             sram_0_avalon_sram_slave_slavearbiterlockenable2;
  wire             sram_0_avalon_sram_slave_unreg_firsttransfer;
  wire             sram_0_avalon_sram_slave_waits_for_read;
  wire             sram_0_avalon_sram_slave_waits_for_write;
  wire             sram_0_avalon_sram_slave_write;
  wire    [ 15: 0] sram_0_avalon_sram_slave_writedata;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock2;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_continuerequest;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_rdv_fifo_output_from_sram_0_avalon_sram_slave;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_saved_grant_sram_0_avalon_sram_slave;
  wire             wait_for_sram_0_avalon_sram_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sram_0_avalon_sram_slave_end_xfer;
    end


  assign sram_0_avalon_sram_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave | cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave | cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave | cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave | cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave | cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave | cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave | video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave));
  //assign sram_0_avalon_sram_slave_readdatavalid_from_sa = sram_0_avalon_sram_slave_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sram_0_avalon_sram_slave_readdatavalid_from_sa = sram_0_avalon_sram_slave_readdatavalid;

  //assign sram_0_avalon_sram_slave_readdata_from_sa = sram_0_avalon_sram_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sram_0_avalon_sram_slave_readdata_from_sa = sram_0_avalon_sram_slave_readdata;

  assign cpu_0_data_master_requests_sram_0_avalon_sram_slave = ({cpu_0_data_master_address_to_slave[24 : 19] , 19'b0} == 25'h1880000) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //sram_0_avalon_sram_slave_arb_share_counter set values, which is an e_mux
  assign sram_0_avalon_sram_slave_arb_share_set_values = (cpu_0_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_0_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_0_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_0_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_0_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_0_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_0_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_0_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave)? 2 :
    (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave)? 2 :
    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave)? 2 :
    1;

  //sram_0_avalon_sram_slave_non_bursting_master_requests mux, which is an e_mux
  assign sram_0_avalon_sram_slave_non_bursting_master_requests = cpu_0_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_2_data_master_requests_sram_0_avalon_sram_slave |
    cpu_2_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_3_data_master_requests_sram_0_avalon_sram_slave |
    cpu_3_instruction_master_requests_sram_0_avalon_sram_slave |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave |
    cpu_0_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_2_data_master_requests_sram_0_avalon_sram_slave |
    cpu_2_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_3_data_master_requests_sram_0_avalon_sram_slave |
    cpu_3_instruction_master_requests_sram_0_avalon_sram_slave |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave |
    cpu_0_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_2_data_master_requests_sram_0_avalon_sram_slave |
    cpu_2_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_3_data_master_requests_sram_0_avalon_sram_slave |
    cpu_3_instruction_master_requests_sram_0_avalon_sram_slave |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave |
    cpu_0_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_2_data_master_requests_sram_0_avalon_sram_slave |
    cpu_2_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_3_data_master_requests_sram_0_avalon_sram_slave |
    cpu_3_instruction_master_requests_sram_0_avalon_sram_slave |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave |
    cpu_0_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_2_data_master_requests_sram_0_avalon_sram_slave |
    cpu_2_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_3_data_master_requests_sram_0_avalon_sram_slave |
    cpu_3_instruction_master_requests_sram_0_avalon_sram_slave |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave |
    cpu_0_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_2_data_master_requests_sram_0_avalon_sram_slave |
    cpu_2_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_3_data_master_requests_sram_0_avalon_sram_slave |
    cpu_3_instruction_master_requests_sram_0_avalon_sram_slave |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave |
    cpu_0_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_2_data_master_requests_sram_0_avalon_sram_slave |
    cpu_2_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_3_data_master_requests_sram_0_avalon_sram_slave |
    cpu_3_instruction_master_requests_sram_0_avalon_sram_slave |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave |
    cpu_0_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_data_master_requests_sram_0_avalon_sram_slave |
    cpu_1_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_2_data_master_requests_sram_0_avalon_sram_slave |
    cpu_2_instruction_master_requests_sram_0_avalon_sram_slave |
    cpu_3_data_master_requests_sram_0_avalon_sram_slave |
    cpu_3_instruction_master_requests_sram_0_avalon_sram_slave |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave;

  //sram_0_avalon_sram_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign sram_0_avalon_sram_slave_any_bursting_master_saved_grant = 0;

  //sram_0_avalon_sram_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign sram_0_avalon_sram_slave_arb_share_counter_next_value = sram_0_avalon_sram_slave_firsttransfer ? (sram_0_avalon_sram_slave_arb_share_set_values - 1) : |sram_0_avalon_sram_slave_arb_share_counter ? (sram_0_avalon_sram_slave_arb_share_counter - 1) : 0;

  //sram_0_avalon_sram_slave_allgrants all slave grants, which is an e_mux
  assign sram_0_avalon_sram_slave_allgrants = (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector) |
    (|sram_0_avalon_sram_slave_grant_vector);

  //sram_0_avalon_sram_slave_end_xfer assignment, which is an e_assign
  assign sram_0_avalon_sram_slave_end_xfer = ~(sram_0_avalon_sram_slave_waits_for_read | sram_0_avalon_sram_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_sram_0_avalon_sram_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_end_xfer & (~sram_0_avalon_sram_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sram_0_avalon_sram_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign sram_0_avalon_sram_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_sram_0_avalon_sram_slave & sram_0_avalon_sram_slave_allgrants) | (end_xfer_arb_share_counter_term_sram_0_avalon_sram_slave & ~sram_0_avalon_sram_slave_non_bursting_master_requests);

  //sram_0_avalon_sram_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sram_0_avalon_sram_slave_arb_share_counter <= 0;
      else if (sram_0_avalon_sram_slave_arb_counter_enable)
          sram_0_avalon_sram_slave_arb_share_counter <= sram_0_avalon_sram_slave_arb_share_counter_next_value;
    end


  //sram_0_avalon_sram_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sram_0_avalon_sram_slave_slavearbiterlockenable <= 0;
      else if ((|sram_0_avalon_sram_slave_master_qreq_vector & end_xfer_arb_share_counter_term_sram_0_avalon_sram_slave) | (end_xfer_arb_share_counter_term_sram_0_avalon_sram_slave & ~sram_0_avalon_sram_slave_non_bursting_master_requests))
          sram_0_avalon_sram_slave_slavearbiterlockenable <= |sram_0_avalon_sram_slave_arb_share_counter_next_value;
    end


  //cpu_0/data_master sram_0/avalon_sram_slave arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = sram_0_avalon_sram_slave_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //sram_0_avalon_sram_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sram_0_avalon_sram_slave_slavearbiterlockenable2 = |sram_0_avalon_sram_slave_arb_share_counter_next_value;

  //cpu_0/data_master sram_0/avalon_sram_slave arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = sram_0_avalon_sram_slave_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_1/data_master sram_0/avalon_sram_slave arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = sram_0_avalon_sram_slave_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master sram_0/avalon_sram_slave arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = sram_0_avalon_sram_slave_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted sram_0/avalon_sram_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_sram_0_avalon_sram_slave <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_sram_0_avalon_sram_slave <= cpu_1_data_master_saved_grant_sram_0_avalon_sram_slave ? 1 : (sram_0_avalon_sram_slave_arbitration_holdoff_internal | ~cpu_1_data_master_requests_sram_0_avalon_sram_slave) ? 0 : last_cycle_cpu_1_data_master_granted_slave_sram_0_avalon_sram_slave;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_data_master_requests_sram_0_avalon_sram_slave);

  //sram_0_avalon_sram_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  assign sram_0_avalon_sram_slave_any_continuerequest = cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_instruction_master_continuerequest |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_1_instruction_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_2_instruction_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_3_instruction_master_continuerequest;

  //cpu_1/instruction_master sram_0/avalon_sram_slave arbiterlock, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock = sram_0_avalon_sram_slave_slavearbiterlockenable & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master sram_0/avalon_sram_slave arbiterlock2, which is an e_assign
  assign cpu_1_instruction_master_arbiterlock2 = sram_0_avalon_sram_slave_slavearbiterlockenable2 & cpu_1_instruction_master_continuerequest;

  //cpu_1/instruction_master granted sram_0/avalon_sram_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_instruction_master_granted_slave_sram_0_avalon_sram_slave <= 0;
      else 
        last_cycle_cpu_1_instruction_master_granted_slave_sram_0_avalon_sram_slave <= cpu_1_instruction_master_saved_grant_sram_0_avalon_sram_slave ? 1 : (sram_0_avalon_sram_slave_arbitration_holdoff_internal | ~cpu_1_instruction_master_requests_sram_0_avalon_sram_slave) ? 0 : last_cycle_cpu_1_instruction_master_granted_slave_sram_0_avalon_sram_slave;
    end


  //cpu_1_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_1_instruction_master_continuerequest = (last_cycle_cpu_1_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_1_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_1_instruction_master_requests_sram_0_avalon_sram_slave);

  //cpu_2/data_master sram_0/avalon_sram_slave arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = sram_0_avalon_sram_slave_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master sram_0/avalon_sram_slave arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = sram_0_avalon_sram_slave_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted sram_0/avalon_sram_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_sram_0_avalon_sram_slave <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_sram_0_avalon_sram_slave <= cpu_2_data_master_saved_grant_sram_0_avalon_sram_slave ? 1 : (sram_0_avalon_sram_slave_arbitration_holdoff_internal | ~cpu_2_data_master_requests_sram_0_avalon_sram_slave) ? 0 : last_cycle_cpu_2_data_master_granted_slave_sram_0_avalon_sram_slave;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_data_master_requests_sram_0_avalon_sram_slave);

  //cpu_2/instruction_master sram_0/avalon_sram_slave arbiterlock, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock = sram_0_avalon_sram_slave_slavearbiterlockenable & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master sram_0/avalon_sram_slave arbiterlock2, which is an e_assign
  assign cpu_2_instruction_master_arbiterlock2 = sram_0_avalon_sram_slave_slavearbiterlockenable2 & cpu_2_instruction_master_continuerequest;

  //cpu_2/instruction_master granted sram_0/avalon_sram_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_instruction_master_granted_slave_sram_0_avalon_sram_slave <= 0;
      else 
        last_cycle_cpu_2_instruction_master_granted_slave_sram_0_avalon_sram_slave <= cpu_2_instruction_master_saved_grant_sram_0_avalon_sram_slave ? 1 : (sram_0_avalon_sram_slave_arbitration_holdoff_internal | ~cpu_2_instruction_master_requests_sram_0_avalon_sram_slave) ? 0 : last_cycle_cpu_2_instruction_master_granted_slave_sram_0_avalon_sram_slave;
    end


  //cpu_2_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_2_instruction_master_continuerequest = (last_cycle_cpu_2_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_2_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_2_instruction_master_requests_sram_0_avalon_sram_slave);

  //cpu_3/data_master sram_0/avalon_sram_slave arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = sram_0_avalon_sram_slave_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master sram_0/avalon_sram_slave arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = sram_0_avalon_sram_slave_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted sram_0/avalon_sram_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_sram_0_avalon_sram_slave <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_sram_0_avalon_sram_slave <= cpu_3_data_master_saved_grant_sram_0_avalon_sram_slave ? 1 : (sram_0_avalon_sram_slave_arbitration_holdoff_internal | ~cpu_3_data_master_requests_sram_0_avalon_sram_slave) ? 0 : last_cycle_cpu_3_data_master_granted_slave_sram_0_avalon_sram_slave;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_data_master_requests_sram_0_avalon_sram_slave);

  //cpu_3/instruction_master sram_0/avalon_sram_slave arbiterlock, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock = sram_0_avalon_sram_slave_slavearbiterlockenable & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master sram_0/avalon_sram_slave arbiterlock2, which is an e_assign
  assign cpu_3_instruction_master_arbiterlock2 = sram_0_avalon_sram_slave_slavearbiterlockenable2 & cpu_3_instruction_master_continuerequest;

  //cpu_3/instruction_master granted sram_0/avalon_sram_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_instruction_master_granted_slave_sram_0_avalon_sram_slave <= 0;
      else 
        last_cycle_cpu_3_instruction_master_granted_slave_sram_0_avalon_sram_slave <= cpu_3_instruction_master_saved_grant_sram_0_avalon_sram_slave ? 1 : (sram_0_avalon_sram_slave_arbitration_holdoff_internal | ~cpu_3_instruction_master_requests_sram_0_avalon_sram_slave) ? 0 : last_cycle_cpu_3_instruction_master_granted_slave_sram_0_avalon_sram_slave;
    end


  //cpu_3_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_3_instruction_master_continuerequest = (last_cycle_cpu_3_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_instruction_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_3_instruction_master_granted_slave_sram_0_avalon_sram_slave & cpu_3_instruction_master_requests_sram_0_avalon_sram_slave);

  //video_pixel_buffer_dma_0/avalon_pixel_dma_master sram_0/avalon_sram_slave arbiterlock2, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock2 = sram_0_avalon_sram_slave_slavearbiterlockenable2 & video_pixel_buffer_dma_0_avalon_pixel_dma_master_continuerequest;

  //video_pixel_buffer_dma_0/avalon_pixel_dma_master granted sram_0/avalon_sram_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_slave_sram_0_avalon_sram_slave <= 0;
      else 
        last_cycle_video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_slave_sram_0_avalon_sram_slave <= video_pixel_buffer_dma_0_avalon_pixel_dma_master_saved_grant_sram_0_avalon_sram_slave ? 1 : (sram_0_avalon_sram_slave_arbitration_holdoff_internal | ~video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave) ? 0 : last_cycle_video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_slave_sram_0_avalon_sram_slave;
    end


  //video_pixel_buffer_dma_0_avalon_pixel_dma_master_continuerequest continued request, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_continuerequest = (last_cycle_video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_slave_sram_0_avalon_sram_slave & video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_slave_sram_0_avalon_sram_slave & video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_slave_sram_0_avalon_sram_slave & video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_slave_sram_0_avalon_sram_slave & video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_slave_sram_0_avalon_sram_slave & video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_slave_sram_0_avalon_sram_slave & video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_slave_sram_0_avalon_sram_slave & video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave);

  assign cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave = cpu_0_data_master_requests_sram_0_avalon_sram_slave & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (1 < cpu_0_data_master_latency_counter))) | ((!cpu_0_data_master_byteenable_sram_0_avalon_sram_slave) & cpu_0_data_master_write) | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock | (video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock & (saved_chosen_master_btw_video_pixel_buffer_dma_0_avalon_pixel_dma_master_and_sram_0_avalon_sram_slave)));
  //unique name for sram_0_avalon_sram_slave_move_on_to_next_transaction, which is an e_assign
  assign sram_0_avalon_sram_slave_move_on_to_next_transaction = sram_0_avalon_sram_slave_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_0_data_master_to_sram_0_avalon_sram_slave, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_0_data_master_to_sram_0_avalon_sram_slave_module rdv_fifo_for_cpu_0_data_master_to_sram_0_avalon_sram_slave
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_0_data_master_granted_sram_0_avalon_sram_slave),
      .data_out             (cpu_0_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave),
      .empty                (),
      .fifo_contains_ones_n (cpu_0_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave),
      .full                 (),
      .read                 (sram_0_avalon_sram_slave_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sram_0_avalon_sram_slave_waits_for_read)
    );

  assign cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register = ~cpu_0_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  //local readdatavalid cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave, which is an e_mux
  assign cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave = (sram_0_avalon_sram_slave_readdatavalid_from_sa & cpu_0_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave) & ~ cpu_0_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;

  //sram_0_avalon_sram_slave_writedata mux, which is an e_mux
  assign sram_0_avalon_sram_slave_writedata = (cpu_0_data_master_granted_sram_0_avalon_sram_slave)? cpu_0_data_master_dbs_write_16 :
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave)? cpu_1_data_master_dbs_write_16 :
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave)? cpu_2_data_master_dbs_write_16 :
    cpu_3_data_master_dbs_write_16;

  assign cpu_1_data_master_requests_sram_0_avalon_sram_slave = ({cpu_1_data_master_address_to_slave[24 : 19] , 19'b0} == 25'h1880000) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //cpu_0/data_master granted sram_0/avalon_sram_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_sram_0_avalon_sram_slave <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_sram_0_avalon_sram_slave <= cpu_0_data_master_saved_grant_sram_0_avalon_sram_slave ? 1 : (sram_0_avalon_sram_slave_arbitration_holdoff_internal | ~cpu_0_data_master_requests_sram_0_avalon_sram_slave) ? 0 : last_cycle_cpu_0_data_master_granted_slave_sram_0_avalon_sram_slave;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_0_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_0_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_0_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_0_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_0_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_0_data_master_requests_sram_0_avalon_sram_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_sram_0_avalon_sram_slave & cpu_0_data_master_requests_sram_0_avalon_sram_slave);

  assign cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave = cpu_1_data_master_requests_sram_0_avalon_sram_slave & ~((cpu_1_data_master_read & ((cpu_1_data_master_latency_counter != 0) | (1 < cpu_1_data_master_latency_counter))) | ((!cpu_1_data_master_byteenable_sram_0_avalon_sram_slave) & cpu_1_data_master_write) | cpu_0_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock | (video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock & (saved_chosen_master_btw_video_pixel_buffer_dma_0_avalon_pixel_dma_master_and_sram_0_avalon_sram_slave)));
  //rdv_fifo_for_cpu_1_data_master_to_sram_0_avalon_sram_slave, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_1_data_master_to_sram_0_avalon_sram_slave_module rdv_fifo_for_cpu_1_data_master_to_sram_0_avalon_sram_slave
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_1_data_master_granted_sram_0_avalon_sram_slave),
      .data_out             (cpu_1_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave),
      .empty                (),
      .fifo_contains_ones_n (cpu_1_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave),
      .full                 (),
      .read                 (sram_0_avalon_sram_slave_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sram_0_avalon_sram_slave_waits_for_read)
    );

  assign cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register = ~cpu_1_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  //local readdatavalid cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave, which is an e_mux
  assign cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave = (sram_0_avalon_sram_slave_readdatavalid_from_sa & cpu_1_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave) & ~ cpu_1_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;

  assign cpu_1_instruction_master_requests_sram_0_avalon_sram_slave = (({cpu_1_instruction_master_address_to_slave[24 : 19] , 19'b0} == 25'h1880000) & (cpu_1_instruction_master_read)) & cpu_1_instruction_master_read;
  assign cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave = cpu_1_instruction_master_requests_sram_0_avalon_sram_slave & ~((cpu_1_instruction_master_read & ((cpu_1_instruction_master_latency_counter != 0) | (1 < cpu_1_instruction_master_latency_counter))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock | (video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock & (saved_chosen_master_btw_video_pixel_buffer_dma_0_avalon_pixel_dma_master_and_sram_0_avalon_sram_slave)));
  //rdv_fifo_for_cpu_1_instruction_master_to_sram_0_avalon_sram_slave, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_1_instruction_master_to_sram_0_avalon_sram_slave_module rdv_fifo_for_cpu_1_instruction_master_to_sram_0_avalon_sram_slave
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave),
      .data_out             (cpu_1_instruction_master_rdv_fifo_output_from_sram_0_avalon_sram_slave),
      .empty                (),
      .fifo_contains_ones_n (cpu_1_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave),
      .full                 (),
      .read                 (sram_0_avalon_sram_slave_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sram_0_avalon_sram_slave_waits_for_read)
    );

  assign cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register = ~cpu_1_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  //local readdatavalid cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave, which is an e_mux
  assign cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave = (sram_0_avalon_sram_slave_readdatavalid_from_sa & cpu_1_instruction_master_rdv_fifo_output_from_sram_0_avalon_sram_slave) & ~ cpu_1_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave;

  assign cpu_2_data_master_requests_sram_0_avalon_sram_slave = ({cpu_2_data_master_address_to_slave[24 : 19] , 19'b0} == 25'h1880000) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave = cpu_2_data_master_requests_sram_0_avalon_sram_slave & ~((cpu_2_data_master_read & ((cpu_2_data_master_latency_counter != 0) | (1 < cpu_2_data_master_latency_counter))) | ((!cpu_2_data_master_byteenable_sram_0_avalon_sram_slave) & cpu_2_data_master_write) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock | (video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock & (saved_chosen_master_btw_video_pixel_buffer_dma_0_avalon_pixel_dma_master_and_sram_0_avalon_sram_slave)));
  //rdv_fifo_for_cpu_2_data_master_to_sram_0_avalon_sram_slave, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_2_data_master_to_sram_0_avalon_sram_slave_module rdv_fifo_for_cpu_2_data_master_to_sram_0_avalon_sram_slave
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_2_data_master_granted_sram_0_avalon_sram_slave),
      .data_out             (cpu_2_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave),
      .empty                (),
      .fifo_contains_ones_n (cpu_2_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave),
      .full                 (),
      .read                 (sram_0_avalon_sram_slave_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sram_0_avalon_sram_slave_waits_for_read)
    );

  assign cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register = ~cpu_2_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  //local readdatavalid cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave, which is an e_mux
  assign cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave = (sram_0_avalon_sram_slave_readdatavalid_from_sa & cpu_2_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave) & ~ cpu_2_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;

  assign cpu_2_instruction_master_requests_sram_0_avalon_sram_slave = (({cpu_2_instruction_master_address_to_slave[24 : 19] , 19'b0} == 25'h1880000) & (cpu_2_instruction_master_read)) & cpu_2_instruction_master_read;
  assign cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave = cpu_2_instruction_master_requests_sram_0_avalon_sram_slave & ~((cpu_2_instruction_master_read & ((cpu_2_instruction_master_latency_counter != 0) | (1 < cpu_2_instruction_master_latency_counter))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock | (video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock & (saved_chosen_master_btw_video_pixel_buffer_dma_0_avalon_pixel_dma_master_and_sram_0_avalon_sram_slave)));
  //rdv_fifo_for_cpu_2_instruction_master_to_sram_0_avalon_sram_slave, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_2_instruction_master_to_sram_0_avalon_sram_slave_module rdv_fifo_for_cpu_2_instruction_master_to_sram_0_avalon_sram_slave
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave),
      .data_out             (cpu_2_instruction_master_rdv_fifo_output_from_sram_0_avalon_sram_slave),
      .empty                (),
      .fifo_contains_ones_n (cpu_2_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave),
      .full                 (),
      .read                 (sram_0_avalon_sram_slave_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sram_0_avalon_sram_slave_waits_for_read)
    );

  assign cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register = ~cpu_2_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  //local readdatavalid cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave, which is an e_mux
  assign cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave = (sram_0_avalon_sram_slave_readdatavalid_from_sa & cpu_2_instruction_master_rdv_fifo_output_from_sram_0_avalon_sram_slave) & ~ cpu_2_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave;

  assign cpu_3_data_master_requests_sram_0_avalon_sram_slave = ({cpu_3_data_master_address_to_slave[24 : 19] , 19'b0} == 25'h1880000) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave = cpu_3_data_master_requests_sram_0_avalon_sram_slave & ~((cpu_3_data_master_read & ((cpu_3_data_master_latency_counter != 0) | (1 < cpu_3_data_master_latency_counter))) | ((!cpu_3_data_master_byteenable_sram_0_avalon_sram_slave) & cpu_3_data_master_write) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_instruction_master_arbiterlock | (video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock & (saved_chosen_master_btw_video_pixel_buffer_dma_0_avalon_pixel_dma_master_and_sram_0_avalon_sram_slave)));
  //rdv_fifo_for_cpu_3_data_master_to_sram_0_avalon_sram_slave, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_3_data_master_to_sram_0_avalon_sram_slave_module rdv_fifo_for_cpu_3_data_master_to_sram_0_avalon_sram_slave
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_3_data_master_granted_sram_0_avalon_sram_slave),
      .data_out             (cpu_3_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave),
      .empty                (),
      .fifo_contains_ones_n (cpu_3_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave),
      .full                 (),
      .read                 (sram_0_avalon_sram_slave_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sram_0_avalon_sram_slave_waits_for_read)
    );

  assign cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register = ~cpu_3_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  //local readdatavalid cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave, which is an e_mux
  assign cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave = (sram_0_avalon_sram_slave_readdatavalid_from_sa & cpu_3_data_master_rdv_fifo_output_from_sram_0_avalon_sram_slave) & ~ cpu_3_data_master_rdv_fifo_empty_sram_0_avalon_sram_slave;

  assign cpu_3_instruction_master_requests_sram_0_avalon_sram_slave = (({cpu_3_instruction_master_address_to_slave[24 : 19] , 19'b0} == 25'h1880000) & (cpu_3_instruction_master_read)) & cpu_3_instruction_master_read;
  assign cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave = cpu_3_instruction_master_requests_sram_0_avalon_sram_slave & ~((cpu_3_instruction_master_read & ((cpu_3_instruction_master_latency_counter != 0) | (1 < cpu_3_instruction_master_latency_counter))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | (video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock & (saved_chosen_master_btw_video_pixel_buffer_dma_0_avalon_pixel_dma_master_and_sram_0_avalon_sram_slave)));
  //rdv_fifo_for_cpu_3_instruction_master_to_sram_0_avalon_sram_slave, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_3_instruction_master_to_sram_0_avalon_sram_slave_module rdv_fifo_for_cpu_3_instruction_master_to_sram_0_avalon_sram_slave
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave),
      .data_out             (cpu_3_instruction_master_rdv_fifo_output_from_sram_0_avalon_sram_slave),
      .empty                (),
      .fifo_contains_ones_n (cpu_3_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave),
      .full                 (),
      .read                 (sram_0_avalon_sram_slave_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sram_0_avalon_sram_slave_waits_for_read)
    );

  assign cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register = ~cpu_3_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  //local readdatavalid cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave, which is an e_mux
  assign cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave = (sram_0_avalon_sram_slave_readdatavalid_from_sa & cpu_3_instruction_master_rdv_fifo_output_from_sram_0_avalon_sram_slave) & ~ cpu_3_instruction_master_rdv_fifo_empty_sram_0_avalon_sram_slave;

  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave = (({video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave[31 : 19] , 19'b0} == 32'h1880000) & (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read)) & video_pixel_buffer_dma_0_avalon_pixel_dma_master_read;
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave = video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave & ~((video_pixel_buffer_dma_0_avalon_pixel_dma_master_read & ((video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter != 0) | (1 < video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_1_instruction_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_2_instruction_master_arbiterlock | cpu_3_data_master_arbiterlock | cpu_3_instruction_master_arbiterlock);
  //rdv_fifo_for_video_pixel_buffer_dma_0_avalon_pixel_dma_master_to_sram_0_avalon_sram_slave, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_video_pixel_buffer_dma_0_avalon_pixel_dma_master_to_sram_0_avalon_sram_slave_module rdv_fifo_for_video_pixel_buffer_dma_0_avalon_pixel_dma_master_to_sram_0_avalon_sram_slave
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave),
      .data_out             (video_pixel_buffer_dma_0_avalon_pixel_dma_master_rdv_fifo_output_from_sram_0_avalon_sram_slave),
      .empty                (),
      .fifo_contains_ones_n (video_pixel_buffer_dma_0_avalon_pixel_dma_master_rdv_fifo_empty_sram_0_avalon_sram_slave),
      .full                 (),
      .read                 (sram_0_avalon_sram_slave_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sram_0_avalon_sram_slave_waits_for_read)
    );

  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave_shift_register = ~video_pixel_buffer_dma_0_avalon_pixel_dma_master_rdv_fifo_empty_sram_0_avalon_sram_slave;
  //local readdatavalid video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave = (sram_0_avalon_sram_slave_readdatavalid_from_sa & video_pixel_buffer_dma_0_avalon_pixel_dma_master_rdv_fifo_output_from_sram_0_avalon_sram_slave) & ~ video_pixel_buffer_dma_0_avalon_pixel_dma_master_rdv_fifo_empty_sram_0_avalon_sram_slave;

  //allow new arb cycle for sram_0/avalon_sram_slave, which is an e_assign
  assign sram_0_avalon_sram_slave_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_1_instruction_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_2_instruction_master_arbiterlock & ~cpu_3_data_master_arbiterlock & ~cpu_3_instruction_master_arbiterlock & ~(video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock & (saved_chosen_master_btw_video_pixel_buffer_dma_0_avalon_pixel_dma_master_and_sram_0_avalon_sram_slave));

  //video_pixel_buffer_dma_0/avalon_pixel_dma_master assignment into master qualified-requests vector for sram_0/avalon_sram_slave, which is an e_assign
  assign sram_0_avalon_sram_slave_master_qreq_vector[0] = video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave;

  //video_pixel_buffer_dma_0/avalon_pixel_dma_master grant sram_0/avalon_sram_slave, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_grant_vector[0];

  //video_pixel_buffer_dma_0/avalon_pixel_dma_master saved-grant sram_0/avalon_sram_slave, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_saved_grant_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_arb_winner[0] && video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave;

  //saved chosen master btw video_pixel_buffer_dma_0/avalon_pixel_dma_master and sram_0/avalon_sram_slave, which is an e_assign
  assign saved_chosen_master_btw_video_pixel_buffer_dma_0_avalon_pixel_dma_master_and_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_saved_chosen_master_vector[0];

  //cpu_3/instruction_master assignment into master qualified-requests vector for sram_0/avalon_sram_slave, which is an e_assign
  assign sram_0_avalon_sram_slave_master_qreq_vector[1] = cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave;

  //cpu_3/instruction_master grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_3_instruction_master_granted_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_grant_vector[1];

  //cpu_3/instruction_master saved-grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_3_instruction_master_saved_grant_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_arb_winner[1] && cpu_3_instruction_master_requests_sram_0_avalon_sram_slave;

  //cpu_3/data_master assignment into master qualified-requests vector for sram_0/avalon_sram_slave, which is an e_assign
  assign sram_0_avalon_sram_slave_master_qreq_vector[2] = cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave;

  //cpu_3/data_master grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_3_data_master_granted_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_grant_vector[2];

  //cpu_3/data_master saved-grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_3_data_master_saved_grant_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_arb_winner[2] && cpu_3_data_master_requests_sram_0_avalon_sram_slave;

  //cpu_2/instruction_master assignment into master qualified-requests vector for sram_0/avalon_sram_slave, which is an e_assign
  assign sram_0_avalon_sram_slave_master_qreq_vector[3] = cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave;

  //cpu_2/instruction_master grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_2_instruction_master_granted_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_grant_vector[3];

  //cpu_2/instruction_master saved-grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_2_instruction_master_saved_grant_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_arb_winner[3] && cpu_2_instruction_master_requests_sram_0_avalon_sram_slave;

  //cpu_2/data_master assignment into master qualified-requests vector for sram_0/avalon_sram_slave, which is an e_assign
  assign sram_0_avalon_sram_slave_master_qreq_vector[4] = cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave;

  //cpu_2/data_master grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_2_data_master_granted_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_grant_vector[4];

  //cpu_2/data_master saved-grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_2_data_master_saved_grant_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_arb_winner[4] && cpu_2_data_master_requests_sram_0_avalon_sram_slave;

  //cpu_1/instruction_master assignment into master qualified-requests vector for sram_0/avalon_sram_slave, which is an e_assign
  assign sram_0_avalon_sram_slave_master_qreq_vector[5] = cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave;

  //cpu_1/instruction_master grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_1_instruction_master_granted_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_grant_vector[5];

  //cpu_1/instruction_master saved-grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_1_instruction_master_saved_grant_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_arb_winner[5] && cpu_1_instruction_master_requests_sram_0_avalon_sram_slave;

  //cpu_1/data_master assignment into master qualified-requests vector for sram_0/avalon_sram_slave, which is an e_assign
  assign sram_0_avalon_sram_slave_master_qreq_vector[6] = cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave;

  //cpu_1/data_master grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_1_data_master_granted_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_grant_vector[6];

  //cpu_1/data_master saved-grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_1_data_master_saved_grant_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_arb_winner[6] && cpu_1_data_master_requests_sram_0_avalon_sram_slave;

  //cpu_0/data_master assignment into master qualified-requests vector for sram_0/avalon_sram_slave, which is an e_assign
  assign sram_0_avalon_sram_slave_master_qreq_vector[7] = cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave;

  //cpu_0/data_master grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_0_data_master_granted_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_grant_vector[7];

  //cpu_0/data_master saved-grant sram_0/avalon_sram_slave, which is an e_assign
  assign cpu_0_data_master_saved_grant_sram_0_avalon_sram_slave = sram_0_avalon_sram_slave_arb_winner[7] && cpu_0_data_master_requests_sram_0_avalon_sram_slave;

  //sram_0/avalon_sram_slave chosen-master double-vector, which is an e_assign
  assign sram_0_avalon_sram_slave_chosen_master_double_vector = {sram_0_avalon_sram_slave_master_qreq_vector, sram_0_avalon_sram_slave_master_qreq_vector} & ({~sram_0_avalon_sram_slave_master_qreq_vector, ~sram_0_avalon_sram_slave_master_qreq_vector} + sram_0_avalon_sram_slave_arb_addend);

  //stable onehot encoding of arb winner
  assign sram_0_avalon_sram_slave_arb_winner = (sram_0_avalon_sram_slave_allow_new_arb_cycle & | sram_0_avalon_sram_slave_grant_vector) ? sram_0_avalon_sram_slave_grant_vector : sram_0_avalon_sram_slave_saved_chosen_master_vector;

  //saved sram_0_avalon_sram_slave_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sram_0_avalon_sram_slave_saved_chosen_master_vector <= 0;
      else if (sram_0_avalon_sram_slave_allow_new_arb_cycle)
          sram_0_avalon_sram_slave_saved_chosen_master_vector <= |sram_0_avalon_sram_slave_grant_vector ? sram_0_avalon_sram_slave_grant_vector : sram_0_avalon_sram_slave_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign sram_0_avalon_sram_slave_grant_vector = {(sram_0_avalon_sram_slave_chosen_master_double_vector[7] | sram_0_avalon_sram_slave_chosen_master_double_vector[15]),
    (sram_0_avalon_sram_slave_chosen_master_double_vector[6] | sram_0_avalon_sram_slave_chosen_master_double_vector[14]),
    (sram_0_avalon_sram_slave_chosen_master_double_vector[5] | sram_0_avalon_sram_slave_chosen_master_double_vector[13]),
    (sram_0_avalon_sram_slave_chosen_master_double_vector[4] | sram_0_avalon_sram_slave_chosen_master_double_vector[12]),
    (sram_0_avalon_sram_slave_chosen_master_double_vector[3] | sram_0_avalon_sram_slave_chosen_master_double_vector[11]),
    (sram_0_avalon_sram_slave_chosen_master_double_vector[2] | sram_0_avalon_sram_slave_chosen_master_double_vector[10]),
    (sram_0_avalon_sram_slave_chosen_master_double_vector[1] | sram_0_avalon_sram_slave_chosen_master_double_vector[9]),
    (sram_0_avalon_sram_slave_chosen_master_double_vector[0] | sram_0_avalon_sram_slave_chosen_master_double_vector[8])};

  //sram_0/avalon_sram_slave chosen master rotated left, which is an e_assign
  assign sram_0_avalon_sram_slave_chosen_master_rot_left = (sram_0_avalon_sram_slave_arb_winner << 1) ? (sram_0_avalon_sram_slave_arb_winner << 1) : 1;

  //sram_0/avalon_sram_slave's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sram_0_avalon_sram_slave_arb_addend <= 1;
      else if (|sram_0_avalon_sram_slave_grant_vector)
          sram_0_avalon_sram_slave_arb_addend <= sram_0_avalon_sram_slave_end_xfer? sram_0_avalon_sram_slave_chosen_master_rot_left : sram_0_avalon_sram_slave_grant_vector;
    end


  //~sram_0_avalon_sram_slave_reset assignment, which is an e_assign
  assign sram_0_avalon_sram_slave_reset = ~reset_n;

  //sram_0_avalon_sram_slave_firsttransfer first transaction, which is an e_assign
  assign sram_0_avalon_sram_slave_firsttransfer = sram_0_avalon_sram_slave_begins_xfer ? sram_0_avalon_sram_slave_unreg_firsttransfer : sram_0_avalon_sram_slave_reg_firsttransfer;

  //sram_0_avalon_sram_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign sram_0_avalon_sram_slave_unreg_firsttransfer = ~(sram_0_avalon_sram_slave_slavearbiterlockenable & sram_0_avalon_sram_slave_any_continuerequest);

  //sram_0_avalon_sram_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sram_0_avalon_sram_slave_reg_firsttransfer <= 1'b1;
      else if (sram_0_avalon_sram_slave_begins_xfer)
          sram_0_avalon_sram_slave_reg_firsttransfer <= sram_0_avalon_sram_slave_unreg_firsttransfer;
    end


  //sram_0_avalon_sram_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sram_0_avalon_sram_slave_beginbursttransfer_internal = sram_0_avalon_sram_slave_begins_xfer;

  //sram_0_avalon_sram_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign sram_0_avalon_sram_slave_arbitration_holdoff_internal = sram_0_avalon_sram_slave_begins_xfer & sram_0_avalon_sram_slave_firsttransfer;

  //sram_0_avalon_sram_slave_read assignment, which is an e_mux
  assign sram_0_avalon_sram_slave_read = (cpu_0_data_master_granted_sram_0_avalon_sram_slave & cpu_0_data_master_read) | (cpu_1_data_master_granted_sram_0_avalon_sram_slave & cpu_1_data_master_read) | (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave & cpu_1_instruction_master_read) | (cpu_2_data_master_granted_sram_0_avalon_sram_slave & cpu_2_data_master_read) | (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave & cpu_2_instruction_master_read) | (cpu_3_data_master_granted_sram_0_avalon_sram_slave & cpu_3_data_master_read) | (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave & cpu_3_instruction_master_read) | (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave & video_pixel_buffer_dma_0_avalon_pixel_dma_master_read);

  //sram_0_avalon_sram_slave_write assignment, which is an e_mux
  assign sram_0_avalon_sram_slave_write = (cpu_0_data_master_granted_sram_0_avalon_sram_slave & cpu_0_data_master_write) | (cpu_1_data_master_granted_sram_0_avalon_sram_slave & cpu_1_data_master_write) | (cpu_2_data_master_granted_sram_0_avalon_sram_slave & cpu_2_data_master_write) | (cpu_3_data_master_granted_sram_0_avalon_sram_slave & cpu_3_data_master_write);

  assign shifted_address_to_sram_0_avalon_sram_slave_from_cpu_0_data_master = {cpu_0_data_master_address_to_slave >> 2,
    cpu_0_data_master_dbs_address[1],
    {1 {1'b0}}};

  //sram_0_avalon_sram_slave_address mux, which is an e_mux
  assign sram_0_avalon_sram_slave_address = (cpu_0_data_master_granted_sram_0_avalon_sram_slave)? (shifted_address_to_sram_0_avalon_sram_slave_from_cpu_0_data_master >> 1) :
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave)? (shifted_address_to_sram_0_avalon_sram_slave_from_cpu_1_data_master >> 1) :
    (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave)? (shifted_address_to_sram_0_avalon_sram_slave_from_cpu_1_instruction_master >> 1) :
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave)? (shifted_address_to_sram_0_avalon_sram_slave_from_cpu_2_data_master >> 1) :
    (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave)? (shifted_address_to_sram_0_avalon_sram_slave_from_cpu_2_instruction_master >> 1) :
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave)? (shifted_address_to_sram_0_avalon_sram_slave_from_cpu_3_data_master >> 1) :
    (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave)? (shifted_address_to_sram_0_avalon_sram_slave_from_cpu_3_instruction_master >> 1) :
    (shifted_address_to_sram_0_avalon_sram_slave_from_video_pixel_buffer_dma_0_avalon_pixel_dma_master >> 1);

  assign shifted_address_to_sram_0_avalon_sram_slave_from_cpu_1_data_master = {cpu_1_data_master_address_to_slave >> 2,
    cpu_1_data_master_dbs_address[1],
    {1 {1'b0}}};

  assign shifted_address_to_sram_0_avalon_sram_slave_from_cpu_1_instruction_master = {cpu_1_instruction_master_address_to_slave >> 2,
    cpu_1_instruction_master_dbs_address[1],
    {1 {1'b0}}};

  assign shifted_address_to_sram_0_avalon_sram_slave_from_cpu_2_data_master = {cpu_2_data_master_address_to_slave >> 2,
    cpu_2_data_master_dbs_address[1],
    {1 {1'b0}}};

  assign shifted_address_to_sram_0_avalon_sram_slave_from_cpu_2_instruction_master = {cpu_2_instruction_master_address_to_slave >> 2,
    cpu_2_instruction_master_dbs_address[1],
    {1 {1'b0}}};

  assign shifted_address_to_sram_0_avalon_sram_slave_from_cpu_3_data_master = {cpu_3_data_master_address_to_slave >> 2,
    cpu_3_data_master_dbs_address[1],
    {1 {1'b0}}};

  assign shifted_address_to_sram_0_avalon_sram_slave_from_cpu_3_instruction_master = {cpu_3_instruction_master_address_to_slave >> 2,
    cpu_3_instruction_master_dbs_address[1],
    {1 {1'b0}}};

  assign shifted_address_to_sram_0_avalon_sram_slave_from_video_pixel_buffer_dma_0_avalon_pixel_dma_master = {video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave >> 2,
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address[1],
    {1 {1'b0}}};

  //d1_sram_0_avalon_sram_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sram_0_avalon_sram_slave_end_xfer <= 1;
      else 
        d1_sram_0_avalon_sram_slave_end_xfer <= sram_0_avalon_sram_slave_end_xfer;
    end


  //sram_0_avalon_sram_slave_waits_for_read in a cycle, which is an e_mux
  assign sram_0_avalon_sram_slave_waits_for_read = sram_0_avalon_sram_slave_in_a_read_cycle & 0;

  //sram_0_avalon_sram_slave_in_a_read_cycle assignment, which is an e_assign
  assign sram_0_avalon_sram_slave_in_a_read_cycle = (cpu_0_data_master_granted_sram_0_avalon_sram_slave & cpu_0_data_master_read) | (cpu_1_data_master_granted_sram_0_avalon_sram_slave & cpu_1_data_master_read) | (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave & cpu_1_instruction_master_read) | (cpu_2_data_master_granted_sram_0_avalon_sram_slave & cpu_2_data_master_read) | (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave & cpu_2_instruction_master_read) | (cpu_3_data_master_granted_sram_0_avalon_sram_slave & cpu_3_data_master_read) | (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave & cpu_3_instruction_master_read) | (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave & video_pixel_buffer_dma_0_avalon_pixel_dma_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sram_0_avalon_sram_slave_in_a_read_cycle;

  //sram_0_avalon_sram_slave_waits_for_write in a cycle, which is an e_mux
  assign sram_0_avalon_sram_slave_waits_for_write = sram_0_avalon_sram_slave_in_a_write_cycle & 0;

  //sram_0_avalon_sram_slave_in_a_write_cycle assignment, which is an e_assign
  assign sram_0_avalon_sram_slave_in_a_write_cycle = (cpu_0_data_master_granted_sram_0_avalon_sram_slave & cpu_0_data_master_write) | (cpu_1_data_master_granted_sram_0_avalon_sram_slave & cpu_1_data_master_write) | (cpu_2_data_master_granted_sram_0_avalon_sram_slave & cpu_2_data_master_write) | (cpu_3_data_master_granted_sram_0_avalon_sram_slave & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sram_0_avalon_sram_slave_in_a_write_cycle;

  assign wait_for_sram_0_avalon_sram_slave_counter = 0;
  //sram_0_avalon_sram_slave_byteenable byte enable port mux, which is an e_mux
  assign sram_0_avalon_sram_slave_byteenable = (cpu_0_data_master_granted_sram_0_avalon_sram_slave)? cpu_0_data_master_byteenable_sram_0_avalon_sram_slave :
    (cpu_1_data_master_granted_sram_0_avalon_sram_slave)? cpu_1_data_master_byteenable_sram_0_avalon_sram_slave :
    (cpu_2_data_master_granted_sram_0_avalon_sram_slave)? cpu_2_data_master_byteenable_sram_0_avalon_sram_slave :
    (cpu_3_data_master_granted_sram_0_avalon_sram_slave)? cpu_3_data_master_byteenable_sram_0_avalon_sram_slave :
    -1;

  assign {cpu_0_data_master_byteenable_sram_0_avalon_sram_slave_segment_1,
cpu_0_data_master_byteenable_sram_0_avalon_sram_slave_segment_0} = cpu_0_data_master_byteenable;
  assign cpu_0_data_master_byteenable_sram_0_avalon_sram_slave = ((cpu_0_data_master_dbs_address[1] == 0))? cpu_0_data_master_byteenable_sram_0_avalon_sram_slave_segment_0 :
    cpu_0_data_master_byteenable_sram_0_avalon_sram_slave_segment_1;

  assign {cpu_1_data_master_byteenable_sram_0_avalon_sram_slave_segment_1,
cpu_1_data_master_byteenable_sram_0_avalon_sram_slave_segment_0} = cpu_1_data_master_byteenable;
  assign cpu_1_data_master_byteenable_sram_0_avalon_sram_slave = ((cpu_1_data_master_dbs_address[1] == 0))? cpu_1_data_master_byteenable_sram_0_avalon_sram_slave_segment_0 :
    cpu_1_data_master_byteenable_sram_0_avalon_sram_slave_segment_1;

  assign {cpu_2_data_master_byteenable_sram_0_avalon_sram_slave_segment_1,
cpu_2_data_master_byteenable_sram_0_avalon_sram_slave_segment_0} = cpu_2_data_master_byteenable;
  assign cpu_2_data_master_byteenable_sram_0_avalon_sram_slave = ((cpu_2_data_master_dbs_address[1] == 0))? cpu_2_data_master_byteenable_sram_0_avalon_sram_slave_segment_0 :
    cpu_2_data_master_byteenable_sram_0_avalon_sram_slave_segment_1;

  assign {cpu_3_data_master_byteenable_sram_0_avalon_sram_slave_segment_1,
cpu_3_data_master_byteenable_sram_0_avalon_sram_slave_segment_0} = cpu_3_data_master_byteenable;
  assign cpu_3_data_master_byteenable_sram_0_avalon_sram_slave = ((cpu_3_data_master_dbs_address[1] == 0))? cpu_3_data_master_byteenable_sram_0_avalon_sram_slave_segment_0 :
    cpu_3_data_master_byteenable_sram_0_avalon_sram_slave_segment_1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sram_0/avalon_sram_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_sram_0_avalon_sram_slave + cpu_1_data_master_granted_sram_0_avalon_sram_slave + cpu_1_instruction_master_granted_sram_0_avalon_sram_slave + cpu_2_data_master_granted_sram_0_avalon_sram_slave + cpu_2_instruction_master_granted_sram_0_avalon_sram_slave + cpu_3_data_master_granted_sram_0_avalon_sram_slave + cpu_3_instruction_master_granted_sram_0_avalon_sram_slave + video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_sram_0_avalon_sram_slave + cpu_1_data_master_saved_grant_sram_0_avalon_sram_slave + cpu_1_instruction_master_saved_grant_sram_0_avalon_sram_slave + cpu_2_data_master_saved_grant_sram_0_avalon_sram_slave + cpu_2_instruction_master_saved_grant_sram_0_avalon_sram_slave + cpu_3_data_master_saved_grant_sram_0_avalon_sram_slave + cpu_3_instruction_master_saved_grant_sram_0_avalon_sram_slave + video_pixel_buffer_dma_0_avalon_pixel_dma_master_saved_grant_sram_0_avalon_sram_slave > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sysid_control_slave_arbitrator (
                                        // inputs:
                                         clk,
                                         cpu_0_data_master_address_to_slave,
                                         cpu_0_data_master_latency_counter,
                                         cpu_0_data_master_read,
                                         cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_0_data_master_write,
                                         cpu_1_data_master_address_to_slave,
                                         cpu_1_data_master_latency_counter,
                                         cpu_1_data_master_read,
                                         cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_1_data_master_write,
                                         cpu_2_data_master_address_to_slave,
                                         cpu_2_data_master_latency_counter,
                                         cpu_2_data_master_read,
                                         cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_2_data_master_write,
                                         cpu_3_data_master_address_to_slave,
                                         cpu_3_data_master_latency_counter,
                                         cpu_3_data_master_read,
                                         cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                         cpu_3_data_master_write,
                                         reset_n,
                                         sysid_control_slave_readdata,

                                        // outputs:
                                         cpu_0_data_master_granted_sysid_control_slave,
                                         cpu_0_data_master_qualified_request_sysid_control_slave,
                                         cpu_0_data_master_read_data_valid_sysid_control_slave,
                                         cpu_0_data_master_requests_sysid_control_slave,
                                         cpu_1_data_master_granted_sysid_control_slave,
                                         cpu_1_data_master_qualified_request_sysid_control_slave,
                                         cpu_1_data_master_read_data_valid_sysid_control_slave,
                                         cpu_1_data_master_requests_sysid_control_slave,
                                         cpu_2_data_master_granted_sysid_control_slave,
                                         cpu_2_data_master_qualified_request_sysid_control_slave,
                                         cpu_2_data_master_read_data_valid_sysid_control_slave,
                                         cpu_2_data_master_requests_sysid_control_slave,
                                         cpu_3_data_master_granted_sysid_control_slave,
                                         cpu_3_data_master_qualified_request_sysid_control_slave,
                                         cpu_3_data_master_read_data_valid_sysid_control_slave,
                                         cpu_3_data_master_requests_sysid_control_slave,
                                         d1_sysid_control_slave_end_xfer,
                                         sysid_control_slave_address,
                                         sysid_control_slave_readdata_from_sa,
                                         sysid_control_slave_reset_n
                                      )
;

  output           cpu_0_data_master_granted_sysid_control_slave;
  output           cpu_0_data_master_qualified_request_sysid_control_slave;
  output           cpu_0_data_master_read_data_valid_sysid_control_slave;
  output           cpu_0_data_master_requests_sysid_control_slave;
  output           cpu_1_data_master_granted_sysid_control_slave;
  output           cpu_1_data_master_qualified_request_sysid_control_slave;
  output           cpu_1_data_master_read_data_valid_sysid_control_slave;
  output           cpu_1_data_master_requests_sysid_control_slave;
  output           cpu_2_data_master_granted_sysid_control_slave;
  output           cpu_2_data_master_qualified_request_sysid_control_slave;
  output           cpu_2_data_master_read_data_valid_sysid_control_slave;
  output           cpu_2_data_master_requests_sysid_control_slave;
  output           cpu_3_data_master_granted_sysid_control_slave;
  output           cpu_3_data_master_qualified_request_sysid_control_slave;
  output           cpu_3_data_master_read_data_valid_sysid_control_slave;
  output           cpu_3_data_master_requests_sysid_control_slave;
  output           d1_sysid_control_slave_end_xfer;
  output           sysid_control_slave_address;
  output  [ 31: 0] sysid_control_slave_readdata_from_sa;
  output           sysid_control_slave_reset_n;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input            reset_n;
  input   [ 31: 0] sysid_control_slave_readdata;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_sysid_control_slave;
  wire             cpu_0_data_master_qualified_request_sysid_control_slave;
  wire             cpu_0_data_master_read_data_valid_sysid_control_slave;
  wire             cpu_0_data_master_requests_sysid_control_slave;
  wire             cpu_0_data_master_saved_grant_sysid_control_slave;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_sysid_control_slave;
  wire             cpu_1_data_master_qualified_request_sysid_control_slave;
  wire             cpu_1_data_master_read_data_valid_sysid_control_slave;
  wire             cpu_1_data_master_requests_sysid_control_slave;
  wire             cpu_1_data_master_saved_grant_sysid_control_slave;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_sysid_control_slave;
  wire             cpu_2_data_master_qualified_request_sysid_control_slave;
  wire             cpu_2_data_master_read_data_valid_sysid_control_slave;
  wire             cpu_2_data_master_requests_sysid_control_slave;
  wire             cpu_2_data_master_saved_grant_sysid_control_slave;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_sysid_control_slave;
  wire             cpu_3_data_master_qualified_request_sysid_control_slave;
  wire             cpu_3_data_master_read_data_valid_sysid_control_slave;
  wire             cpu_3_data_master_requests_sysid_control_slave;
  wire             cpu_3_data_master_saved_grant_sysid_control_slave;
  reg              d1_reasons_to_wait;
  reg              d1_sysid_control_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sysid_control_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_sysid_control_slave;
  reg              last_cycle_cpu_1_data_master_granted_slave_sysid_control_slave;
  reg              last_cycle_cpu_2_data_master_granted_slave_sysid_control_slave;
  reg              last_cycle_cpu_3_data_master_granted_slave_sysid_control_slave;
  wire    [ 24: 0] shifted_address_to_sysid_control_slave_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_sysid_control_slave_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_sysid_control_slave_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_sysid_control_slave_from_cpu_3_data_master;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_allgrants;
  wire             sysid_control_slave_allow_new_arb_cycle;
  wire             sysid_control_slave_any_bursting_master_saved_grant;
  wire             sysid_control_slave_any_continuerequest;
  reg     [  3: 0] sysid_control_slave_arb_addend;
  wire             sysid_control_slave_arb_counter_enable;
  reg     [  2: 0] sysid_control_slave_arb_share_counter;
  wire    [  2: 0] sysid_control_slave_arb_share_counter_next_value;
  wire    [  2: 0] sysid_control_slave_arb_share_set_values;
  wire    [  3: 0] sysid_control_slave_arb_winner;
  wire             sysid_control_slave_arbitration_holdoff_internal;
  wire             sysid_control_slave_beginbursttransfer_internal;
  wire             sysid_control_slave_begins_xfer;
  wire    [  7: 0] sysid_control_slave_chosen_master_double_vector;
  wire    [  3: 0] sysid_control_slave_chosen_master_rot_left;
  wire             sysid_control_slave_end_xfer;
  wire             sysid_control_slave_firsttransfer;
  wire    [  3: 0] sysid_control_slave_grant_vector;
  wire             sysid_control_slave_in_a_read_cycle;
  wire             sysid_control_slave_in_a_write_cycle;
  wire    [  3: 0] sysid_control_slave_master_qreq_vector;
  wire             sysid_control_slave_non_bursting_master_requests;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  reg              sysid_control_slave_reg_firsttransfer;
  wire             sysid_control_slave_reset_n;
  reg     [  3: 0] sysid_control_slave_saved_chosen_master_vector;
  reg              sysid_control_slave_slavearbiterlockenable;
  wire             sysid_control_slave_slavearbiterlockenable2;
  wire             sysid_control_slave_unreg_firsttransfer;
  wire             sysid_control_slave_waits_for_read;
  wire             sysid_control_slave_waits_for_write;
  wire             wait_for_sysid_control_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sysid_control_slave_end_xfer;
    end


  assign sysid_control_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_sysid_control_slave | cpu_1_data_master_qualified_request_sysid_control_slave | cpu_2_data_master_qualified_request_sysid_control_slave | cpu_3_data_master_qualified_request_sysid_control_slave));
  //assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata;

  assign cpu_0_data_master_requests_sysid_control_slave = (({cpu_0_data_master_address_to_slave[24 : 3] , 3'b0} == 25'h19030c0) & (cpu_0_data_master_read | cpu_0_data_master_write)) & cpu_0_data_master_read;
  //sysid_control_slave_arb_share_counter set values, which is an e_mux
  assign sysid_control_slave_arb_share_set_values = 1;

  //sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  assign sysid_control_slave_non_bursting_master_requests = cpu_0_data_master_requests_sysid_control_slave |
    cpu_1_data_master_requests_sysid_control_slave |
    cpu_2_data_master_requests_sysid_control_slave |
    cpu_3_data_master_requests_sysid_control_slave |
    cpu_0_data_master_requests_sysid_control_slave |
    cpu_1_data_master_requests_sysid_control_slave |
    cpu_2_data_master_requests_sysid_control_slave |
    cpu_3_data_master_requests_sysid_control_slave |
    cpu_0_data_master_requests_sysid_control_slave |
    cpu_1_data_master_requests_sysid_control_slave |
    cpu_2_data_master_requests_sysid_control_slave |
    cpu_3_data_master_requests_sysid_control_slave |
    cpu_0_data_master_requests_sysid_control_slave |
    cpu_1_data_master_requests_sysid_control_slave |
    cpu_2_data_master_requests_sysid_control_slave |
    cpu_3_data_master_requests_sysid_control_slave;

  //sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign sysid_control_slave_any_bursting_master_saved_grant = 0;

  //sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign sysid_control_slave_arb_share_counter_next_value = sysid_control_slave_firsttransfer ? (sysid_control_slave_arb_share_set_values - 1) : |sysid_control_slave_arb_share_counter ? (sysid_control_slave_arb_share_counter - 1) : 0;

  //sysid_control_slave_allgrants all slave grants, which is an e_mux
  assign sysid_control_slave_allgrants = (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector) |
    (|sysid_control_slave_grant_vector);

  //sysid_control_slave_end_xfer assignment, which is an e_assign
  assign sysid_control_slave_end_xfer = ~(sysid_control_slave_waits_for_read | sysid_control_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sysid_control_slave = sysid_control_slave_end_xfer & (~sysid_control_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign sysid_control_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_sysid_control_slave & sysid_control_slave_allgrants) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests);

  //sysid_control_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_arb_share_counter <= 0;
      else if (sysid_control_slave_arb_counter_enable)
          sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
    end


  //sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_slavearbiterlockenable <= 0;
      else if ((|sysid_control_slave_master_qreq_vector & end_xfer_arb_share_counter_term_sysid_control_slave) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests))
          sysid_control_slave_slavearbiterlockenable <= |sysid_control_slave_arb_share_counter_next_value;
    end


  //cpu_0/data_master sysid/control_slave arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = sysid_control_slave_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sysid_control_slave_slavearbiterlockenable2 = |sysid_control_slave_arb_share_counter_next_value;

  //cpu_0/data_master sysid/control_slave arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = sysid_control_slave_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_1/data_master sysid/control_slave arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = sysid_control_slave_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master sysid/control_slave arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = sysid_control_slave_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted sysid/control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_sysid_control_slave <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_sysid_control_slave <= cpu_1_data_master_saved_grant_sysid_control_slave ? 1 : (sysid_control_slave_arbitration_holdoff_internal | ~cpu_1_data_master_requests_sysid_control_slave) ? 0 : last_cycle_cpu_1_data_master_granted_slave_sysid_control_slave;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_sysid_control_slave & cpu_1_data_master_requests_sysid_control_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_sysid_control_slave & cpu_1_data_master_requests_sysid_control_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_sysid_control_slave & cpu_1_data_master_requests_sysid_control_slave);

  //sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  assign sysid_control_slave_any_continuerequest = cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest;

  //cpu_2/data_master sysid/control_slave arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = sysid_control_slave_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master sysid/control_slave arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = sysid_control_slave_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted sysid/control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_sysid_control_slave <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_sysid_control_slave <= cpu_2_data_master_saved_grant_sysid_control_slave ? 1 : (sysid_control_slave_arbitration_holdoff_internal | ~cpu_2_data_master_requests_sysid_control_slave) ? 0 : last_cycle_cpu_2_data_master_granted_slave_sysid_control_slave;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_sysid_control_slave & cpu_2_data_master_requests_sysid_control_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_sysid_control_slave & cpu_2_data_master_requests_sysid_control_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_sysid_control_slave & cpu_2_data_master_requests_sysid_control_slave);

  //cpu_3/data_master sysid/control_slave arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = sysid_control_slave_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master sysid/control_slave arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = sysid_control_slave_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted sysid/control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_sysid_control_slave <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_sysid_control_slave <= cpu_3_data_master_saved_grant_sysid_control_slave ? 1 : (sysid_control_slave_arbitration_holdoff_internal | ~cpu_3_data_master_requests_sysid_control_slave) ? 0 : last_cycle_cpu_3_data_master_granted_slave_sysid_control_slave;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_sysid_control_slave & cpu_3_data_master_requests_sysid_control_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_sysid_control_slave & cpu_3_data_master_requests_sysid_control_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_sysid_control_slave & cpu_3_data_master_requests_sysid_control_slave);

  assign cpu_0_data_master_qualified_request_sysid_control_slave = cpu_0_data_master_requests_sysid_control_slave & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_sysid_control_slave, which is an e_mux
  assign cpu_0_data_master_read_data_valid_sysid_control_slave = cpu_0_data_master_granted_sysid_control_slave & cpu_0_data_master_read & ~sysid_control_slave_waits_for_read;

  assign cpu_1_data_master_requests_sysid_control_slave = (({cpu_1_data_master_address_to_slave[24 : 3] , 3'b0} == 25'h19030c0) & (cpu_1_data_master_read | cpu_1_data_master_write)) & cpu_1_data_master_read;
  //cpu_0/data_master granted sysid/control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_sysid_control_slave <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_sysid_control_slave <= cpu_0_data_master_saved_grant_sysid_control_slave ? 1 : (sysid_control_slave_arbitration_holdoff_internal | ~cpu_0_data_master_requests_sysid_control_slave) ? 0 : last_cycle_cpu_0_data_master_granted_slave_sysid_control_slave;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_sysid_control_slave & cpu_0_data_master_requests_sysid_control_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_sysid_control_slave & cpu_0_data_master_requests_sysid_control_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_sysid_control_slave & cpu_0_data_master_requests_sysid_control_slave);

  assign cpu_1_data_master_qualified_request_sysid_control_slave = cpu_1_data_master_requests_sysid_control_slave & ~((cpu_1_data_master_read & ((cpu_1_data_master_latency_counter != 0) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_1_data_master_read_data_valid_sysid_control_slave, which is an e_mux
  assign cpu_1_data_master_read_data_valid_sysid_control_slave = cpu_1_data_master_granted_sysid_control_slave & cpu_1_data_master_read & ~sysid_control_slave_waits_for_read;

  assign cpu_2_data_master_requests_sysid_control_slave = (({cpu_2_data_master_address_to_slave[24 : 3] , 3'b0} == 25'h19030c0) & (cpu_2_data_master_read | cpu_2_data_master_write)) & cpu_2_data_master_read;
  assign cpu_2_data_master_qualified_request_sysid_control_slave = cpu_2_data_master_requests_sysid_control_slave & ~((cpu_2_data_master_read & ((cpu_2_data_master_latency_counter != 0) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //local readdatavalid cpu_2_data_master_read_data_valid_sysid_control_slave, which is an e_mux
  assign cpu_2_data_master_read_data_valid_sysid_control_slave = cpu_2_data_master_granted_sysid_control_slave & cpu_2_data_master_read & ~sysid_control_slave_waits_for_read;

  assign cpu_3_data_master_requests_sysid_control_slave = (({cpu_3_data_master_address_to_slave[24 : 3] , 3'b0} == 25'h19030c0) & (cpu_3_data_master_read | cpu_3_data_master_write)) & cpu_3_data_master_read;
  assign cpu_3_data_master_qualified_request_sysid_control_slave = cpu_3_data_master_requests_sysid_control_slave & ~((cpu_3_data_master_read & ((cpu_3_data_master_latency_counter != 0) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock);
  //local readdatavalid cpu_3_data_master_read_data_valid_sysid_control_slave, which is an e_mux
  assign cpu_3_data_master_read_data_valid_sysid_control_slave = cpu_3_data_master_granted_sysid_control_slave & cpu_3_data_master_read & ~sysid_control_slave_waits_for_read;

  //allow new arb cycle for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_3_data_master_arbiterlock;

  //cpu_3/data_master assignment into master qualified-requests vector for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_master_qreq_vector[0] = cpu_3_data_master_qualified_request_sysid_control_slave;

  //cpu_3/data_master grant sysid/control_slave, which is an e_assign
  assign cpu_3_data_master_granted_sysid_control_slave = sysid_control_slave_grant_vector[0];

  //cpu_3/data_master saved-grant sysid/control_slave, which is an e_assign
  assign cpu_3_data_master_saved_grant_sysid_control_slave = sysid_control_slave_arb_winner[0] && cpu_3_data_master_requests_sysid_control_slave;

  //cpu_2/data_master assignment into master qualified-requests vector for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_master_qreq_vector[1] = cpu_2_data_master_qualified_request_sysid_control_slave;

  //cpu_2/data_master grant sysid/control_slave, which is an e_assign
  assign cpu_2_data_master_granted_sysid_control_slave = sysid_control_slave_grant_vector[1];

  //cpu_2/data_master saved-grant sysid/control_slave, which is an e_assign
  assign cpu_2_data_master_saved_grant_sysid_control_slave = sysid_control_slave_arb_winner[1] && cpu_2_data_master_requests_sysid_control_slave;

  //cpu_1/data_master assignment into master qualified-requests vector for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_master_qreq_vector[2] = cpu_1_data_master_qualified_request_sysid_control_slave;

  //cpu_1/data_master grant sysid/control_slave, which is an e_assign
  assign cpu_1_data_master_granted_sysid_control_slave = sysid_control_slave_grant_vector[2];

  //cpu_1/data_master saved-grant sysid/control_slave, which is an e_assign
  assign cpu_1_data_master_saved_grant_sysid_control_slave = sysid_control_slave_arb_winner[2] && cpu_1_data_master_requests_sysid_control_slave;

  //cpu_0/data_master assignment into master qualified-requests vector for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_master_qreq_vector[3] = cpu_0_data_master_qualified_request_sysid_control_slave;

  //cpu_0/data_master grant sysid/control_slave, which is an e_assign
  assign cpu_0_data_master_granted_sysid_control_slave = sysid_control_slave_grant_vector[3];

  //cpu_0/data_master saved-grant sysid/control_slave, which is an e_assign
  assign cpu_0_data_master_saved_grant_sysid_control_slave = sysid_control_slave_arb_winner[3] && cpu_0_data_master_requests_sysid_control_slave;

  //sysid/control_slave chosen-master double-vector, which is an e_assign
  assign sysid_control_slave_chosen_master_double_vector = {sysid_control_slave_master_qreq_vector, sysid_control_slave_master_qreq_vector} & ({~sysid_control_slave_master_qreq_vector, ~sysid_control_slave_master_qreq_vector} + sysid_control_slave_arb_addend);

  //stable onehot encoding of arb winner
  assign sysid_control_slave_arb_winner = (sysid_control_slave_allow_new_arb_cycle & | sysid_control_slave_grant_vector) ? sysid_control_slave_grant_vector : sysid_control_slave_saved_chosen_master_vector;

  //saved sysid_control_slave_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_saved_chosen_master_vector <= 0;
      else if (sysid_control_slave_allow_new_arb_cycle)
          sysid_control_slave_saved_chosen_master_vector <= |sysid_control_slave_grant_vector ? sysid_control_slave_grant_vector : sysid_control_slave_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign sysid_control_slave_grant_vector = {(sysid_control_slave_chosen_master_double_vector[3] | sysid_control_slave_chosen_master_double_vector[7]),
    (sysid_control_slave_chosen_master_double_vector[2] | sysid_control_slave_chosen_master_double_vector[6]),
    (sysid_control_slave_chosen_master_double_vector[1] | sysid_control_slave_chosen_master_double_vector[5]),
    (sysid_control_slave_chosen_master_double_vector[0] | sysid_control_slave_chosen_master_double_vector[4])};

  //sysid/control_slave chosen master rotated left, which is an e_assign
  assign sysid_control_slave_chosen_master_rot_left = (sysid_control_slave_arb_winner << 1) ? (sysid_control_slave_arb_winner << 1) : 1;

  //sysid/control_slave's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_arb_addend <= 1;
      else if (|sysid_control_slave_grant_vector)
          sysid_control_slave_arb_addend <= sysid_control_slave_end_xfer? sysid_control_slave_chosen_master_rot_left : sysid_control_slave_grant_vector;
    end


  //sysid_control_slave_reset_n assignment, which is an e_assign
  assign sysid_control_slave_reset_n = reset_n;

  //sysid_control_slave_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_firsttransfer = sysid_control_slave_begins_xfer ? sysid_control_slave_unreg_firsttransfer : sysid_control_slave_reg_firsttransfer;

  //sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_unreg_firsttransfer = ~(sysid_control_slave_slavearbiterlockenable & sysid_control_slave_any_continuerequest);

  //sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_reg_firsttransfer <= 1'b1;
      else if (sysid_control_slave_begins_xfer)
          sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
    end


  //sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sysid_control_slave_beginbursttransfer_internal = sysid_control_slave_begins_xfer;

  //sysid_control_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign sysid_control_slave_arbitration_holdoff_internal = sysid_control_slave_begins_xfer & sysid_control_slave_firsttransfer;

  assign shifted_address_to_sysid_control_slave_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //sysid_control_slave_address mux, which is an e_mux
  assign sysid_control_slave_address = (cpu_0_data_master_granted_sysid_control_slave)? (shifted_address_to_sysid_control_slave_from_cpu_0_data_master >> 2) :
    (cpu_1_data_master_granted_sysid_control_slave)? (shifted_address_to_sysid_control_slave_from_cpu_1_data_master >> 2) :
    (cpu_2_data_master_granted_sysid_control_slave)? (shifted_address_to_sysid_control_slave_from_cpu_2_data_master >> 2) :
    (shifted_address_to_sysid_control_slave_from_cpu_3_data_master >> 2);

  assign shifted_address_to_sysid_control_slave_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_sysid_control_slave_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_sysid_control_slave_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  //d1_sysid_control_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sysid_control_slave_end_xfer <= 1;
      else 
        d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end


  //sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_read = sysid_control_slave_in_a_read_cycle & sysid_control_slave_begins_xfer;

  //sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_read_cycle = (cpu_0_data_master_granted_sysid_control_slave & cpu_0_data_master_read) | (cpu_1_data_master_granted_sysid_control_slave & cpu_1_data_master_read) | (cpu_2_data_master_granted_sysid_control_slave & cpu_2_data_master_read) | (cpu_3_data_master_granted_sysid_control_slave & cpu_3_data_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sysid_control_slave_in_a_read_cycle;

  //sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_write = sysid_control_slave_in_a_write_cycle & 0;

  //sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_write_cycle = (cpu_0_data_master_granted_sysid_control_slave & cpu_0_data_master_write) | (cpu_1_data_master_granted_sysid_control_slave & cpu_1_data_master_write) | (cpu_2_data_master_granted_sysid_control_slave & cpu_2_data_master_write) | (cpu_3_data_master_granted_sysid_control_slave & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sysid_control_slave_in_a_write_cycle;

  assign wait_for_sysid_control_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sysid/control_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_sysid_control_slave + cpu_1_data_master_granted_sysid_control_slave + cpu_2_data_master_granted_sysid_control_slave + cpu_3_data_master_granted_sysid_control_slave > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_sysid_control_slave + cpu_1_data_master_saved_grant_sysid_control_slave + cpu_2_data_master_saved_grant_sysid_control_slave + cpu_3_data_master_saved_grant_sysid_control_slave > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module video_dual_clock_buffer_0_avalon_dc_buffer_sink_arbitrator (
                                                                    // inputs:
                                                                     clk,
                                                                     reset_n,
                                                                     video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready,
                                                                     video_scaler_0_avalon_scaler_source_data,
                                                                     video_scaler_0_avalon_scaler_source_endofpacket,
                                                                     video_scaler_0_avalon_scaler_source_startofpacket,
                                                                     video_scaler_0_avalon_scaler_source_valid,

                                                                    // outputs:
                                                                     video_dual_clock_buffer_0_avalon_dc_buffer_sink_data,
                                                                     video_dual_clock_buffer_0_avalon_dc_buffer_sink_endofpacket,
                                                                     video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa,
                                                                     video_dual_clock_buffer_0_avalon_dc_buffer_sink_startofpacket,
                                                                     video_dual_clock_buffer_0_avalon_dc_buffer_sink_valid
                                                                  )
;

  output  [ 29: 0] video_dual_clock_buffer_0_avalon_dc_buffer_sink_data;
  output           video_dual_clock_buffer_0_avalon_dc_buffer_sink_endofpacket;
  output           video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa;
  output           video_dual_clock_buffer_0_avalon_dc_buffer_sink_startofpacket;
  output           video_dual_clock_buffer_0_avalon_dc_buffer_sink_valid;
  input            clk;
  input            reset_n;
  input            video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready;
  input   [ 29: 0] video_scaler_0_avalon_scaler_source_data;
  input            video_scaler_0_avalon_scaler_source_endofpacket;
  input            video_scaler_0_avalon_scaler_source_startofpacket;
  input            video_scaler_0_avalon_scaler_source_valid;

  wire    [ 29: 0] video_dual_clock_buffer_0_avalon_dc_buffer_sink_data;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_sink_endofpacket;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_sink_startofpacket;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_sink_valid;
  //mux video_dual_clock_buffer_0_avalon_dc_buffer_sink_data, which is an e_mux
  assign video_dual_clock_buffer_0_avalon_dc_buffer_sink_data = video_scaler_0_avalon_scaler_source_data;

  //mux video_dual_clock_buffer_0_avalon_dc_buffer_sink_endofpacket, which is an e_mux
  assign video_dual_clock_buffer_0_avalon_dc_buffer_sink_endofpacket = video_scaler_0_avalon_scaler_source_endofpacket;

  //assign video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa = video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa = video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready;

  //mux video_dual_clock_buffer_0_avalon_dc_buffer_sink_startofpacket, which is an e_mux
  assign video_dual_clock_buffer_0_avalon_dc_buffer_sink_startofpacket = video_scaler_0_avalon_scaler_source_startofpacket;

  //mux video_dual_clock_buffer_0_avalon_dc_buffer_sink_valid, which is an e_mux
  assign video_dual_clock_buffer_0_avalon_dc_buffer_sink_valid = video_scaler_0_avalon_scaler_source_valid;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module video_dual_clock_buffer_0_avalon_dc_buffer_source_arbitrator (
                                                                      // inputs:
                                                                       clk,
                                                                       reset_n,
                                                                       video_dual_clock_buffer_0_avalon_dc_buffer_source_data,
                                                                       video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket,
                                                                       video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket,
                                                                       video_dual_clock_buffer_0_avalon_dc_buffer_source_valid,
                                                                       video_vga_controller_0_avalon_vga_sink_ready_from_sa,

                                                                      // outputs:
                                                                       video_dual_clock_buffer_0_avalon_dc_buffer_source_ready
                                                                    )
;

  output           video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;
  input            clk;
  input            reset_n;
  input   [ 29: 0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;
  input            video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;
  input            video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;
  input            video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;
  input            video_vga_controller_0_avalon_vga_sink_ready_from_sa;

  wire             video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;
  //mux video_dual_clock_buffer_0_avalon_dc_buffer_source_ready, which is an e_mux
  assign video_dual_clock_buffer_0_avalon_dc_buffer_source_ready = video_vga_controller_0_avalon_vga_sink_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module video_pixel_buffer_dma_0_avalon_control_slave_arbitrator (
                                                                  // inputs:
                                                                   clk,
                                                                   cpu_0_data_master_address_to_slave,
                                                                   cpu_0_data_master_byteenable,
                                                                   cpu_0_data_master_latency_counter,
                                                                   cpu_0_data_master_read,
                                                                   cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                                   cpu_0_data_master_write,
                                                                   cpu_0_data_master_writedata,
                                                                   cpu_1_data_master_address_to_slave,
                                                                   cpu_1_data_master_byteenable,
                                                                   cpu_1_data_master_latency_counter,
                                                                   cpu_1_data_master_read,
                                                                   cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                                   cpu_1_data_master_write,
                                                                   cpu_1_data_master_writedata,
                                                                   cpu_2_data_master_address_to_slave,
                                                                   cpu_2_data_master_byteenable,
                                                                   cpu_2_data_master_latency_counter,
                                                                   cpu_2_data_master_read,
                                                                   cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                                   cpu_2_data_master_write,
                                                                   cpu_2_data_master_writedata,
                                                                   cpu_3_data_master_address_to_slave,
                                                                   cpu_3_data_master_byteenable,
                                                                   cpu_3_data_master_latency_counter,
                                                                   cpu_3_data_master_read,
                                                                   cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                                   cpu_3_data_master_write,
                                                                   cpu_3_data_master_writedata,
                                                                   reset_n,
                                                                   video_pixel_buffer_dma_0_avalon_control_slave_readdata,

                                                                  // outputs:
                                                                   cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave,
                                                                   d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer,
                                                                   video_pixel_buffer_dma_0_avalon_control_slave_address,
                                                                   video_pixel_buffer_dma_0_avalon_control_slave_byteenable,
                                                                   video_pixel_buffer_dma_0_avalon_control_slave_read,
                                                                   video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa,
                                                                   video_pixel_buffer_dma_0_avalon_control_slave_write,
                                                                   video_pixel_buffer_dma_0_avalon_control_slave_writedata
                                                                )
;

  output           cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  output           cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  output           d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer;
  output  [  1: 0] video_pixel_buffer_dma_0_avalon_control_slave_address;
  output  [  3: 0] video_pixel_buffer_dma_0_avalon_control_slave_byteenable;
  output           video_pixel_buffer_dma_0_avalon_control_slave_read;
  output  [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa;
  output           video_pixel_buffer_dma_0_avalon_control_slave_write;
  output  [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input            cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_1_data_master_address_to_slave;
  input   [  3: 0] cpu_1_data_master_byteenable;
  input            cpu_1_data_master_latency_counter;
  input            cpu_1_data_master_read;
  input            cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_1_data_master_write;
  input   [ 31: 0] cpu_1_data_master_writedata;
  input   [ 24: 0] cpu_2_data_master_address_to_slave;
  input   [  3: 0] cpu_2_data_master_byteenable;
  input            cpu_2_data_master_latency_counter;
  input            cpu_2_data_master_read;
  input            cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_2_data_master_write;
  input   [ 31: 0] cpu_2_data_master_writedata;
  input   [ 24: 0] cpu_3_data_master_address_to_slave;
  input   [  3: 0] cpu_3_data_master_byteenable;
  input            cpu_3_data_master_latency_counter;
  input            cpu_3_data_master_read;
  input            cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            cpu_3_data_master_write;
  input   [ 31: 0] cpu_3_data_master_writedata;
  input            reset_n;
  input   [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_readdata;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  reg              cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
  wire             cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in;
  wire             cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_0_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_1_data_master_arbiterlock;
  wire             cpu_1_data_master_arbiterlock2;
  wire             cpu_1_data_master_continuerequest;
  wire             cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  reg              cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
  wire             cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in;
  wire             cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_1_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_2_data_master_arbiterlock;
  wire             cpu_2_data_master_arbiterlock2;
  wire             cpu_2_data_master_continuerequest;
  wire             cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  reg              cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
  wire             cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in;
  wire             cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_2_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_3_data_master_arbiterlock;
  wire             cpu_3_data_master_arbiterlock2;
  wire             cpu_3_data_master_continuerequest;
  wire             cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  reg              cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
  wire             cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in;
  wire             cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_3_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave;
  reg              d1_reasons_to_wait;
  reg              d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave;
  reg              last_cycle_cpu_1_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave;
  reg              last_cycle_cpu_2_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave;
  reg              last_cycle_cpu_3_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             p1_cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
  wire             p1_cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
  wire             p1_cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
  wire             p1_cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
  wire    [ 24: 0] shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_1_data_master;
  wire    [ 24: 0] shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_2_data_master;
  wire    [ 24: 0] shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_3_data_master;
  wire    [  1: 0] video_pixel_buffer_dma_0_avalon_control_slave_address;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_allgrants;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_allow_new_arb_cycle;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_any_bursting_master_saved_grant;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_any_continuerequest;
  reg     [  3: 0] video_pixel_buffer_dma_0_avalon_control_slave_arb_addend;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_arb_counter_enable;
  reg     [  2: 0] video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter;
  wire    [  2: 0] video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter_next_value;
  wire    [  2: 0] video_pixel_buffer_dma_0_avalon_control_slave_arb_share_set_values;
  wire    [  3: 0] video_pixel_buffer_dma_0_avalon_control_slave_arb_winner;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_arbitration_holdoff_internal;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_beginbursttransfer_internal;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_begins_xfer;
  wire    [  3: 0] video_pixel_buffer_dma_0_avalon_control_slave_byteenable;
  wire    [  7: 0] video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_double_vector;
  wire    [  3: 0] video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_rot_left;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_end_xfer;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_firsttransfer;
  wire    [  3: 0] video_pixel_buffer_dma_0_avalon_control_slave_grant_vector;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_in_a_read_cycle;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_in_a_write_cycle;
  wire    [  3: 0] video_pixel_buffer_dma_0_avalon_control_slave_master_qreq_vector;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_non_bursting_master_requests;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_read;
  wire    [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa;
  reg              video_pixel_buffer_dma_0_avalon_control_slave_reg_firsttransfer;
  reg     [  3: 0] video_pixel_buffer_dma_0_avalon_control_slave_saved_chosen_master_vector;
  reg              video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable2;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_unreg_firsttransfer;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_waits_for_read;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_waits_for_write;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_write;
  wire    [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_writedata;
  wire             wait_for_video_pixel_buffer_dma_0_avalon_control_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~video_pixel_buffer_dma_0_avalon_control_slave_end_xfer;
    end


  assign video_pixel_buffer_dma_0_avalon_control_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave | cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave));
  //assign video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa = video_pixel_buffer_dma_0_avalon_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa = video_pixel_buffer_dma_0_avalon_control_slave_readdata;

  assign cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h19030b0) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter set values, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_arb_share_set_values = 1;

  //video_pixel_buffer_dma_0_avalon_control_slave_non_bursting_master_requests mux, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_non_bursting_master_requests = cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave |
    cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;

  //video_pixel_buffer_dma_0_avalon_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_any_bursting_master_saved_grant = 0;

  //video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter_next_value = video_pixel_buffer_dma_0_avalon_control_slave_firsttransfer ? (video_pixel_buffer_dma_0_avalon_control_slave_arb_share_set_values - 1) : |video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter ? (video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter - 1) : 0;

  //video_pixel_buffer_dma_0_avalon_control_slave_allgrants all slave grants, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_allgrants = (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) |
    (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector);

  //video_pixel_buffer_dma_0_avalon_control_slave_end_xfer assignment, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_end_xfer = ~(video_pixel_buffer_dma_0_avalon_control_slave_waits_for_read | video_pixel_buffer_dma_0_avalon_control_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_video_pixel_buffer_dma_0_avalon_control_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_video_pixel_buffer_dma_0_avalon_control_slave = video_pixel_buffer_dma_0_avalon_control_slave_end_xfer & (~video_pixel_buffer_dma_0_avalon_control_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_video_pixel_buffer_dma_0_avalon_control_slave & video_pixel_buffer_dma_0_avalon_control_slave_allgrants) | (end_xfer_arb_share_counter_term_video_pixel_buffer_dma_0_avalon_control_slave & ~video_pixel_buffer_dma_0_avalon_control_slave_non_bursting_master_requests);

  //video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter <= 0;
      else if (video_pixel_buffer_dma_0_avalon_control_slave_arb_counter_enable)
          video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter <= video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter_next_value;
    end


  //video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable <= 0;
      else if ((|video_pixel_buffer_dma_0_avalon_control_slave_master_qreq_vector & end_xfer_arb_share_counter_term_video_pixel_buffer_dma_0_avalon_control_slave) | (end_xfer_arb_share_counter_term_video_pixel_buffer_dma_0_avalon_control_slave & ~video_pixel_buffer_dma_0_avalon_control_slave_non_bursting_master_requests))
          video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable <= |video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter_next_value;
    end


  //cpu_0/data_master video_pixel_buffer_dma_0/avalon_control_slave arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable2 = |video_pixel_buffer_dma_0_avalon_control_slave_arb_share_counter_next_value;

  //cpu_0/data_master video_pixel_buffer_dma_0/avalon_control_slave arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_1/data_master video_pixel_buffer_dma_0/avalon_control_slave arbiterlock, which is an e_assign
  assign cpu_1_data_master_arbiterlock = video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable & cpu_1_data_master_continuerequest;

  //cpu_1/data_master video_pixel_buffer_dma_0/avalon_control_slave arbiterlock2, which is an e_assign
  assign cpu_1_data_master_arbiterlock2 = video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable2 & cpu_1_data_master_continuerequest;

  //cpu_1/data_master granted video_pixel_buffer_dma_0/avalon_control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_1_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave <= 0;
      else 
        last_cycle_cpu_1_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave <= cpu_1_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave ? 1 : (video_pixel_buffer_dma_0_avalon_control_slave_arbitration_holdoff_internal | ~cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) ? 0 : last_cycle_cpu_1_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave;
    end


  //cpu_1_data_master_continuerequest continued request, which is an e_mux
  assign cpu_1_data_master_continuerequest = (last_cycle_cpu_1_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) |
    (last_cycle_cpu_1_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave);

  //video_pixel_buffer_dma_0_avalon_control_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_any_continuerequest = cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_2_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_3_data_master_continuerequest |
    cpu_0_data_master_continuerequest |
    cpu_1_data_master_continuerequest |
    cpu_2_data_master_continuerequest;

  //cpu_2/data_master video_pixel_buffer_dma_0/avalon_control_slave arbiterlock, which is an e_assign
  assign cpu_2_data_master_arbiterlock = video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable & cpu_2_data_master_continuerequest;

  //cpu_2/data_master video_pixel_buffer_dma_0/avalon_control_slave arbiterlock2, which is an e_assign
  assign cpu_2_data_master_arbiterlock2 = video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable2 & cpu_2_data_master_continuerequest;

  //cpu_2/data_master granted video_pixel_buffer_dma_0/avalon_control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_2_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave <= 0;
      else 
        last_cycle_cpu_2_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave <= cpu_2_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave ? 1 : (video_pixel_buffer_dma_0_avalon_control_slave_arbitration_holdoff_internal | ~cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) ? 0 : last_cycle_cpu_2_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave;
    end


  //cpu_2_data_master_continuerequest continued request, which is an e_mux
  assign cpu_2_data_master_continuerequest = (last_cycle_cpu_2_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) |
    (last_cycle_cpu_2_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave);

  //cpu_3/data_master video_pixel_buffer_dma_0/avalon_control_slave arbiterlock, which is an e_assign
  assign cpu_3_data_master_arbiterlock = video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable & cpu_3_data_master_continuerequest;

  //cpu_3/data_master video_pixel_buffer_dma_0/avalon_control_slave arbiterlock2, which is an e_assign
  assign cpu_3_data_master_arbiterlock2 = video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable2 & cpu_3_data_master_continuerequest;

  //cpu_3/data_master granted video_pixel_buffer_dma_0/avalon_control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_3_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave <= 0;
      else 
        last_cycle_cpu_3_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave <= cpu_3_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave ? 1 : (video_pixel_buffer_dma_0_avalon_control_slave_arbitration_holdoff_internal | ~cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) ? 0 : last_cycle_cpu_3_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave;
    end


  //cpu_3_data_master_continuerequest continued request, which is an e_mux
  assign cpu_3_data_master_continuerequest = (last_cycle_cpu_3_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) |
    (last_cycle_cpu_3_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave);

  assign cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave = cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave & ~((cpu_0_data_master_read & ((1 < cpu_0_data_master_latency_counter) | (|cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in = cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_0_data_master_read & ~video_pixel_buffer_dma_0_avalon_control_slave_waits_for_read;

  //shift register p1 cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register = {cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register, cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in};

  //cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register <= 0;
      else 
        cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register <= p1_cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
    end


  //local readdatavalid cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave, which is an e_mux
  assign cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave = cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;

  //video_pixel_buffer_dma_0_avalon_control_slave_writedata mux, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_writedata = (cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave)? cpu_0_data_master_writedata :
    (cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave)? cpu_1_data_master_writedata :
    (cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave)? cpu_2_data_master_writedata :
    cpu_3_data_master_writedata;

  assign cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave = ({cpu_1_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h19030b0) & (cpu_1_data_master_read | cpu_1_data_master_write);
  //cpu_0/data_master granted video_pixel_buffer_dma_0/avalon_control_slave last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave <= cpu_0_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave ? 1 : (video_pixel_buffer_dma_0_avalon_control_slave_arbitration_holdoff_internal | ~cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) ? 0 : last_cycle_cpu_0_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = (last_cycle_cpu_0_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave) |
    (last_cycle_cpu_0_data_master_granted_slave_video_pixel_buffer_dma_0_avalon_control_slave & cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave);

  assign cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave = cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave & ~((cpu_1_data_master_read & ((1 < cpu_1_data_master_latency_counter) | (|cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_2_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in = cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_1_data_master_read & ~video_pixel_buffer_dma_0_avalon_control_slave_waits_for_read;

  //shift register p1 cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register = {cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register, cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in};

  //cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register <= 0;
      else 
        cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register <= p1_cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
    end


  //local readdatavalid cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave, which is an e_mux
  assign cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave = cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;

  assign cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave = ({cpu_2_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h19030b0) & (cpu_2_data_master_read | cpu_2_data_master_write);
  assign cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave = cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave & ~((cpu_2_data_master_read & ((1 < cpu_2_data_master_latency_counter) | (|cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_3_data_master_arbiterlock);
  //cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in = cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_2_data_master_read & ~video_pixel_buffer_dma_0_avalon_control_slave_waits_for_read;

  //shift register p1 cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register = {cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register, cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in};

  //cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register <= 0;
      else 
        cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register <= p1_cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
    end


  //local readdatavalid cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave, which is an e_mux
  assign cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave = cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;

  assign cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave = ({cpu_3_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h19030b0) & (cpu_3_data_master_read | cpu_3_data_master_write);
  assign cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave = cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave & ~((cpu_3_data_master_read & ((1 < cpu_3_data_master_latency_counter) | (|cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register))) | cpu_0_data_master_arbiterlock | cpu_1_data_master_arbiterlock | cpu_2_data_master_arbiterlock);
  //cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in = cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_3_data_master_read & ~video_pixel_buffer_dma_0_avalon_control_slave_waits_for_read;

  //shift register p1 cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register = {cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register, cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register_in};

  //cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register <= 0;
      else 
        cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register <= p1_cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;
    end


  //local readdatavalid cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave, which is an e_mux
  assign cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave = cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave_shift_register;

  //allow new arb cycle for video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_1_data_master_arbiterlock & ~cpu_2_data_master_arbiterlock & ~cpu_3_data_master_arbiterlock;

  //cpu_3/data_master assignment into master qualified-requests vector for video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_master_qreq_vector[0] = cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;

  //cpu_3/data_master grant video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave = video_pixel_buffer_dma_0_avalon_control_slave_grant_vector[0];

  //cpu_3/data_master saved-grant video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign cpu_3_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave = video_pixel_buffer_dma_0_avalon_control_slave_arb_winner[0] && cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;

  //cpu_2/data_master assignment into master qualified-requests vector for video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_master_qreq_vector[1] = cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;

  //cpu_2/data_master grant video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave = video_pixel_buffer_dma_0_avalon_control_slave_grant_vector[1];

  //cpu_2/data_master saved-grant video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign cpu_2_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave = video_pixel_buffer_dma_0_avalon_control_slave_arb_winner[1] && cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;

  //cpu_1/data_master assignment into master qualified-requests vector for video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_master_qreq_vector[2] = cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;

  //cpu_1/data_master grant video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave = video_pixel_buffer_dma_0_avalon_control_slave_grant_vector[2];

  //cpu_1/data_master saved-grant video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign cpu_1_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave = video_pixel_buffer_dma_0_avalon_control_slave_arb_winner[2] && cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;

  //cpu_0/data_master assignment into master qualified-requests vector for video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_master_qreq_vector[3] = cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;

  //cpu_0/data_master grant video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave = video_pixel_buffer_dma_0_avalon_control_slave_grant_vector[3];

  //cpu_0/data_master saved-grant video_pixel_buffer_dma_0/avalon_control_slave, which is an e_assign
  assign cpu_0_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave = video_pixel_buffer_dma_0_avalon_control_slave_arb_winner[3] && cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;

  //video_pixel_buffer_dma_0/avalon_control_slave chosen-master double-vector, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_double_vector = {video_pixel_buffer_dma_0_avalon_control_slave_master_qreq_vector, video_pixel_buffer_dma_0_avalon_control_slave_master_qreq_vector} & ({~video_pixel_buffer_dma_0_avalon_control_slave_master_qreq_vector, ~video_pixel_buffer_dma_0_avalon_control_slave_master_qreq_vector} + video_pixel_buffer_dma_0_avalon_control_slave_arb_addend);

  //stable onehot encoding of arb winner
  assign video_pixel_buffer_dma_0_avalon_control_slave_arb_winner = (video_pixel_buffer_dma_0_avalon_control_slave_allow_new_arb_cycle & | video_pixel_buffer_dma_0_avalon_control_slave_grant_vector) ? video_pixel_buffer_dma_0_avalon_control_slave_grant_vector : video_pixel_buffer_dma_0_avalon_control_slave_saved_chosen_master_vector;

  //saved video_pixel_buffer_dma_0_avalon_control_slave_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          video_pixel_buffer_dma_0_avalon_control_slave_saved_chosen_master_vector <= 0;
      else if (video_pixel_buffer_dma_0_avalon_control_slave_allow_new_arb_cycle)
          video_pixel_buffer_dma_0_avalon_control_slave_saved_chosen_master_vector <= |video_pixel_buffer_dma_0_avalon_control_slave_grant_vector ? video_pixel_buffer_dma_0_avalon_control_slave_grant_vector : video_pixel_buffer_dma_0_avalon_control_slave_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign video_pixel_buffer_dma_0_avalon_control_slave_grant_vector = {(video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_double_vector[3] | video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_double_vector[7]),
    (video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_double_vector[2] | video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_double_vector[6]),
    (video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_double_vector[1] | video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_double_vector[5]),
    (video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_double_vector[0] | video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_double_vector[4])};

  //video_pixel_buffer_dma_0/avalon_control_slave chosen master rotated left, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_rot_left = (video_pixel_buffer_dma_0_avalon_control_slave_arb_winner << 1) ? (video_pixel_buffer_dma_0_avalon_control_slave_arb_winner << 1) : 1;

  //video_pixel_buffer_dma_0/avalon_control_slave's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          video_pixel_buffer_dma_0_avalon_control_slave_arb_addend <= 1;
      else if (|video_pixel_buffer_dma_0_avalon_control_slave_grant_vector)
          video_pixel_buffer_dma_0_avalon_control_slave_arb_addend <= video_pixel_buffer_dma_0_avalon_control_slave_end_xfer? video_pixel_buffer_dma_0_avalon_control_slave_chosen_master_rot_left : video_pixel_buffer_dma_0_avalon_control_slave_grant_vector;
    end


  //video_pixel_buffer_dma_0_avalon_control_slave_firsttransfer first transaction, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_firsttransfer = video_pixel_buffer_dma_0_avalon_control_slave_begins_xfer ? video_pixel_buffer_dma_0_avalon_control_slave_unreg_firsttransfer : video_pixel_buffer_dma_0_avalon_control_slave_reg_firsttransfer;

  //video_pixel_buffer_dma_0_avalon_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_unreg_firsttransfer = ~(video_pixel_buffer_dma_0_avalon_control_slave_slavearbiterlockenable & video_pixel_buffer_dma_0_avalon_control_slave_any_continuerequest);

  //video_pixel_buffer_dma_0_avalon_control_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          video_pixel_buffer_dma_0_avalon_control_slave_reg_firsttransfer <= 1'b1;
      else if (video_pixel_buffer_dma_0_avalon_control_slave_begins_xfer)
          video_pixel_buffer_dma_0_avalon_control_slave_reg_firsttransfer <= video_pixel_buffer_dma_0_avalon_control_slave_unreg_firsttransfer;
    end


  //video_pixel_buffer_dma_0_avalon_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_beginbursttransfer_internal = video_pixel_buffer_dma_0_avalon_control_slave_begins_xfer;

  //video_pixel_buffer_dma_0_avalon_control_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_arbitration_holdoff_internal = video_pixel_buffer_dma_0_avalon_control_slave_begins_xfer & video_pixel_buffer_dma_0_avalon_control_slave_firsttransfer;

  //video_pixel_buffer_dma_0_avalon_control_slave_read assignment, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_read = (cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_0_data_master_read) | (cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_1_data_master_read) | (cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_2_data_master_read) | (cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_3_data_master_read);

  //video_pixel_buffer_dma_0_avalon_control_slave_write assignment, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_write = (cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_0_data_master_write) | (cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_1_data_master_write) | (cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_2_data_master_write) | (cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_3_data_master_write);

  assign shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //video_pixel_buffer_dma_0_avalon_control_slave_address mux, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_address = (cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave)? (shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_0_data_master >> 2) :
    (cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave)? (shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_1_data_master >> 2) :
    (cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave)? (shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_2_data_master >> 2) :
    (shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_3_data_master >> 2);

  assign shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_1_data_master = cpu_1_data_master_address_to_slave;
  assign shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_2_data_master = cpu_2_data_master_address_to_slave;
  assign shifted_address_to_video_pixel_buffer_dma_0_avalon_control_slave_from_cpu_3_data_master = cpu_3_data_master_address_to_slave;
  //d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer <= 1;
      else 
        d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer <= video_pixel_buffer_dma_0_avalon_control_slave_end_xfer;
    end


  //video_pixel_buffer_dma_0_avalon_control_slave_waits_for_read in a cycle, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_waits_for_read = video_pixel_buffer_dma_0_avalon_control_slave_in_a_read_cycle & 0;

  //video_pixel_buffer_dma_0_avalon_control_slave_in_a_read_cycle assignment, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_in_a_read_cycle = (cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_0_data_master_read) | (cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_1_data_master_read) | (cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_2_data_master_read) | (cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_3_data_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = video_pixel_buffer_dma_0_avalon_control_slave_in_a_read_cycle;

  //video_pixel_buffer_dma_0_avalon_control_slave_waits_for_write in a cycle, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_waits_for_write = video_pixel_buffer_dma_0_avalon_control_slave_in_a_write_cycle & 0;

  //video_pixel_buffer_dma_0_avalon_control_slave_in_a_write_cycle assignment, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_control_slave_in_a_write_cycle = (cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_0_data_master_write) | (cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_1_data_master_write) | (cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_2_data_master_write) | (cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave & cpu_3_data_master_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = video_pixel_buffer_dma_0_avalon_control_slave_in_a_write_cycle;

  assign wait_for_video_pixel_buffer_dma_0_avalon_control_slave_counter = 0;
  //video_pixel_buffer_dma_0_avalon_control_slave_byteenable byte enable port mux, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_control_slave_byteenable = (cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave)? cpu_0_data_master_byteenable :
    (cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave)? cpu_1_data_master_byteenable :
    (cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave)? cpu_2_data_master_byteenable :
    (cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave)? cpu_3_data_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //video_pixel_buffer_dma_0/avalon_control_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave + cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave + cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave + cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave + cpu_1_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave + cpu_2_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave + cpu_3_data_master_saved_grant_video_pixel_buffer_dma_0_avalon_control_slave > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbitrator (
                                                                     // inputs:
                                                                      clk,
                                                                      d1_sram_0_avalon_sram_slave_end_xfer,
                                                                      reset_n,
                                                                      sram_0_avalon_sram_slave_readdata_from_sa,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_address,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_read,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave_shift_register,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave,

                                                                     // outputs:
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_reset,
                                                                      video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest
                                                                   )
;

  output  [ 31: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave;
  output  [  1: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address;
  output           video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter;
  output  [ 31: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata;
  output           video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid;
  output           video_pixel_buffer_dma_0_avalon_pixel_dma_master_reset;
  output           video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest;
  input            clk;
  input            d1_sram_0_avalon_sram_slave_end_xfer;
  input            reset_n;
  input   [ 15: 0] sram_0_avalon_sram_slave_readdata_from_sa;
  input   [ 31: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address;
  input            video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave;
  input            video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave;
  input            video_pixel_buffer_dma_0_avalon_pixel_dma_master_read;
  input            video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave;
  input            video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  input            video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave;

  reg              active_and_waiting_last_time;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire             latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             p1_video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter;
  wire             pre_dbs_count_enable;
  wire             pre_flush_video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid;
  wire             r_3;
  reg     [ 31: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_last_time;
  wire    [ 31: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave;
  reg     [  1: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address;
  wire    [  1: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_increment;
  reg     [  1: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_rdv_counter;
  wire    [  1: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_rdv_counter_inc;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_is_granted_some_slave;
  reg              video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter;
  wire    [  1: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_next_dbs_rdv_counter;
  reg              video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_but_no_slave_selected;
  reg              video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_last_time;
  wire    [ 31: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_reset;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_run;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest;
  //r_3 master_run cascaded wait assignment, which is an e_assign
  assign r_3 = 1 & (video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave | ~video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave) & (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave | ~video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave) & ((~video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave | ~video_pixel_buffer_dma_0_avalon_pixel_dma_master_read | (1 & (video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address[1]) & video_pixel_buffer_dma_0_avalon_pixel_dma_master_read)));

  //cascaded wait assignment, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_run = r_3;

  //optimize select-logic by passing only those address bits which matter.
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave = {13'b110001,
    video_pixel_buffer_dma_0_avalon_pixel_dma_master_address[18 : 0]};

  //video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_but_no_slave_selected <= 0;
      else 
        video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_but_no_slave_selected <= video_pixel_buffer_dma_0_avalon_pixel_dma_master_read & video_pixel_buffer_dma_0_avalon_pixel_dma_master_run & ~video_pixel_buffer_dma_0_avalon_pixel_dma_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_is_granted_some_slave = video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid = video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave & dbs_rdv_counter_overflow;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid = video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_but_no_slave_selected |
    pre_flush_video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid;

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = sram_0_avalon_sram_slave_readdata_from_sa;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //video_pixel_buffer_dma_0/avalon_pixel_dma_master readdata mux, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata = {sram_0_avalon_sram_slave_readdata_from_sa[15 : 0],
    dbs_latent_16_reg_segment_0};

  //actual waitrequest port, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest = ~video_pixel_buffer_dma_0_avalon_pixel_dma_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter <= 0;
      else 
        video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter <= p1_video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter = ((video_pixel_buffer_dma_0_avalon_pixel_dma_master_run & video_pixel_buffer_dma_0_avalon_pixel_dma_master_read))? latency_load_value :
    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter)? video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //~video_pixel_buffer_dma_0_avalon_pixel_dma_master_reset assignment, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_reset = ~reset_n;

  //dbs count increment, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_increment = (video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address + video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address <= 0;
      else if (dbs_count_enable)
          video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address <= next_dbs_address;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_next_dbs_rdv_counter = video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_rdv_counter + video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_rdv_counter_inc;

  //video_pixel_buffer_dma_0_avalon_pixel_dma_master_rdv_inc_mux, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_rdv_counter_inc = 2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_rdv_counter <= video_pixel_buffer_dma_0_avalon_pixel_dma_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_rdv_counter[1] & ~video_pixel_buffer_dma_0_avalon_pixel_dma_master_next_dbs_rdv_counter[1];

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave & video_pixel_buffer_dma_0_avalon_pixel_dma_master_read & 1 & 1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //video_pixel_buffer_dma_0_avalon_pixel_dma_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_last_time <= 0;
      else 
        video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_last_time <= video_pixel_buffer_dma_0_avalon_pixel_dma_master_address;
    end


  //video_pixel_buffer_dma_0/avalon_pixel_dma_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest & (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read);
    end


  //video_pixel_buffer_dma_0_avalon_pixel_dma_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address != video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_last_time))
        begin
          $write("%0d ns: video_pixel_buffer_dma_0_avalon_pixel_dma_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //video_pixel_buffer_dma_0_avalon_pixel_dma_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_last_time <= 0;
      else 
        video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_last_time <= video_pixel_buffer_dma_0_avalon_pixel_dma_master_read;
    end


  //video_pixel_buffer_dma_0_avalon_pixel_dma_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read != video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_last_time))
        begin
          $write("%0d ns: video_pixel_buffer_dma_0_avalon_pixel_dma_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module video_pixel_buffer_dma_0_avalon_pixel_source_arbitrator (
                                                                 // inputs:
                                                                  clk,
                                                                  reset_n,
                                                                  video_pixel_buffer_dma_0_avalon_pixel_source_data,
                                                                  video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket,
                                                                  video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket,
                                                                  video_pixel_buffer_dma_0_avalon_pixel_source_valid,
                                                                  video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa,

                                                                 // outputs:
                                                                  video_pixel_buffer_dma_0_avalon_pixel_source_ready
                                                               )
;

  output           video_pixel_buffer_dma_0_avalon_pixel_source_ready;
  input            clk;
  input            reset_n;
  input   [ 23: 0] video_pixel_buffer_dma_0_avalon_pixel_source_data;
  input            video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket;
  input            video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket;
  input            video_pixel_buffer_dma_0_avalon_pixel_source_valid;
  input            video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa;

  wire             video_pixel_buffer_dma_0_avalon_pixel_source_ready;
  //mux video_pixel_buffer_dma_0_avalon_pixel_source_ready, which is an e_mux
  assign video_pixel_buffer_dma_0_avalon_pixel_source_ready = video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module video_rgb_resampler_0_avalon_rgb_sink_arbitrator (
                                                          // inputs:
                                                           clk,
                                                           reset_n,
                                                           video_pixel_buffer_dma_0_avalon_pixel_source_data,
                                                           video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket,
                                                           video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket,
                                                           video_pixel_buffer_dma_0_avalon_pixel_source_valid,
                                                           video_rgb_resampler_0_avalon_rgb_sink_ready,

                                                          // outputs:
                                                           video_rgb_resampler_0_avalon_rgb_sink_data,
                                                           video_rgb_resampler_0_avalon_rgb_sink_endofpacket,
                                                           video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa,
                                                           video_rgb_resampler_0_avalon_rgb_sink_reset,
                                                           video_rgb_resampler_0_avalon_rgb_sink_startofpacket,
                                                           video_rgb_resampler_0_avalon_rgb_sink_valid
                                                        )
;

  output  [ 23: 0] video_rgb_resampler_0_avalon_rgb_sink_data;
  output           video_rgb_resampler_0_avalon_rgb_sink_endofpacket;
  output           video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa;
  output           video_rgb_resampler_0_avalon_rgb_sink_reset;
  output           video_rgb_resampler_0_avalon_rgb_sink_startofpacket;
  output           video_rgb_resampler_0_avalon_rgb_sink_valid;
  input            clk;
  input            reset_n;
  input   [ 23: 0] video_pixel_buffer_dma_0_avalon_pixel_source_data;
  input            video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket;
  input            video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket;
  input            video_pixel_buffer_dma_0_avalon_pixel_source_valid;
  input            video_rgb_resampler_0_avalon_rgb_sink_ready;

  wire    [ 23: 0] video_rgb_resampler_0_avalon_rgb_sink_data;
  wire             video_rgb_resampler_0_avalon_rgb_sink_endofpacket;
  wire             video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa;
  wire             video_rgb_resampler_0_avalon_rgb_sink_reset;
  wire             video_rgb_resampler_0_avalon_rgb_sink_startofpacket;
  wire             video_rgb_resampler_0_avalon_rgb_sink_valid;
  //mux video_rgb_resampler_0_avalon_rgb_sink_data, which is an e_mux
  assign video_rgb_resampler_0_avalon_rgb_sink_data = video_pixel_buffer_dma_0_avalon_pixel_source_data;

  //mux video_rgb_resampler_0_avalon_rgb_sink_endofpacket, which is an e_mux
  assign video_rgb_resampler_0_avalon_rgb_sink_endofpacket = video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket;

  //assign video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa = video_rgb_resampler_0_avalon_rgb_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa = video_rgb_resampler_0_avalon_rgb_sink_ready;

  //mux video_rgb_resampler_0_avalon_rgb_sink_startofpacket, which is an e_mux
  assign video_rgb_resampler_0_avalon_rgb_sink_startofpacket = video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket;

  //mux video_rgb_resampler_0_avalon_rgb_sink_valid, which is an e_mux
  assign video_rgb_resampler_0_avalon_rgb_sink_valid = video_pixel_buffer_dma_0_avalon_pixel_source_valid;

  //~video_rgb_resampler_0_avalon_rgb_sink_reset assignment, which is an e_assign
  assign video_rgb_resampler_0_avalon_rgb_sink_reset = ~reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module video_rgb_resampler_0_avalon_rgb_source_arbitrator (
                                                            // inputs:
                                                             clk,
                                                             reset_n,
                                                             video_rgb_resampler_0_avalon_rgb_source_data,
                                                             video_rgb_resampler_0_avalon_rgb_source_endofpacket,
                                                             video_rgb_resampler_0_avalon_rgb_source_startofpacket,
                                                             video_rgb_resampler_0_avalon_rgb_source_valid,
                                                             video_scaler_0_avalon_scaler_sink_ready_from_sa,

                                                            // outputs:
                                                             video_rgb_resampler_0_avalon_rgb_source_ready
                                                          )
;

  output           video_rgb_resampler_0_avalon_rgb_source_ready;
  input            clk;
  input            reset_n;
  input   [ 29: 0] video_rgb_resampler_0_avalon_rgb_source_data;
  input            video_rgb_resampler_0_avalon_rgb_source_endofpacket;
  input            video_rgb_resampler_0_avalon_rgb_source_startofpacket;
  input            video_rgb_resampler_0_avalon_rgb_source_valid;
  input            video_scaler_0_avalon_scaler_sink_ready_from_sa;

  wire             video_rgb_resampler_0_avalon_rgb_source_ready;
  //mux video_rgb_resampler_0_avalon_rgb_source_ready, which is an e_mux
  assign video_rgb_resampler_0_avalon_rgb_source_ready = video_scaler_0_avalon_scaler_sink_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module video_scaler_0_avalon_scaler_sink_arbitrator (
                                                      // inputs:
                                                       clk,
                                                       reset_n,
                                                       video_rgb_resampler_0_avalon_rgb_source_data,
                                                       video_rgb_resampler_0_avalon_rgb_source_endofpacket,
                                                       video_rgb_resampler_0_avalon_rgb_source_startofpacket,
                                                       video_rgb_resampler_0_avalon_rgb_source_valid,
                                                       video_scaler_0_avalon_scaler_sink_ready,

                                                      // outputs:
                                                       video_scaler_0_avalon_scaler_sink_data,
                                                       video_scaler_0_avalon_scaler_sink_endofpacket,
                                                       video_scaler_0_avalon_scaler_sink_ready_from_sa,
                                                       video_scaler_0_avalon_scaler_sink_reset,
                                                       video_scaler_0_avalon_scaler_sink_startofpacket,
                                                       video_scaler_0_avalon_scaler_sink_valid
                                                    )
;

  output  [ 29: 0] video_scaler_0_avalon_scaler_sink_data;
  output           video_scaler_0_avalon_scaler_sink_endofpacket;
  output           video_scaler_0_avalon_scaler_sink_ready_from_sa;
  output           video_scaler_0_avalon_scaler_sink_reset;
  output           video_scaler_0_avalon_scaler_sink_startofpacket;
  output           video_scaler_0_avalon_scaler_sink_valid;
  input            clk;
  input            reset_n;
  input   [ 29: 0] video_rgb_resampler_0_avalon_rgb_source_data;
  input            video_rgb_resampler_0_avalon_rgb_source_endofpacket;
  input            video_rgb_resampler_0_avalon_rgb_source_startofpacket;
  input            video_rgb_resampler_0_avalon_rgb_source_valid;
  input            video_scaler_0_avalon_scaler_sink_ready;

  wire    [ 29: 0] video_scaler_0_avalon_scaler_sink_data;
  wire             video_scaler_0_avalon_scaler_sink_endofpacket;
  wire             video_scaler_0_avalon_scaler_sink_ready_from_sa;
  wire             video_scaler_0_avalon_scaler_sink_reset;
  wire             video_scaler_0_avalon_scaler_sink_startofpacket;
  wire             video_scaler_0_avalon_scaler_sink_valid;
  //mux video_scaler_0_avalon_scaler_sink_data, which is an e_mux
  assign video_scaler_0_avalon_scaler_sink_data = video_rgb_resampler_0_avalon_rgb_source_data;

  //mux video_scaler_0_avalon_scaler_sink_endofpacket, which is an e_mux
  assign video_scaler_0_avalon_scaler_sink_endofpacket = video_rgb_resampler_0_avalon_rgb_source_endofpacket;

  //assign video_scaler_0_avalon_scaler_sink_ready_from_sa = video_scaler_0_avalon_scaler_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign video_scaler_0_avalon_scaler_sink_ready_from_sa = video_scaler_0_avalon_scaler_sink_ready;

  //mux video_scaler_0_avalon_scaler_sink_startofpacket, which is an e_mux
  assign video_scaler_0_avalon_scaler_sink_startofpacket = video_rgb_resampler_0_avalon_rgb_source_startofpacket;

  //mux video_scaler_0_avalon_scaler_sink_valid, which is an e_mux
  assign video_scaler_0_avalon_scaler_sink_valid = video_rgb_resampler_0_avalon_rgb_source_valid;

  //~video_scaler_0_avalon_scaler_sink_reset assignment, which is an e_assign
  assign video_scaler_0_avalon_scaler_sink_reset = ~reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module video_scaler_0_avalon_scaler_source_arbitrator (
                                                        // inputs:
                                                         clk,
                                                         reset_n,
                                                         video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa,
                                                         video_scaler_0_avalon_scaler_source_data,
                                                         video_scaler_0_avalon_scaler_source_endofpacket,
                                                         video_scaler_0_avalon_scaler_source_startofpacket,
                                                         video_scaler_0_avalon_scaler_source_valid,

                                                        // outputs:
                                                         video_scaler_0_avalon_scaler_source_ready
                                                      )
;

  output           video_scaler_0_avalon_scaler_source_ready;
  input            clk;
  input            reset_n;
  input            video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa;
  input   [ 29: 0] video_scaler_0_avalon_scaler_source_data;
  input            video_scaler_0_avalon_scaler_source_endofpacket;
  input            video_scaler_0_avalon_scaler_source_startofpacket;
  input            video_scaler_0_avalon_scaler_source_valid;

  wire             video_scaler_0_avalon_scaler_source_ready;
  //mux video_scaler_0_avalon_scaler_source_ready, which is an e_mux
  assign video_scaler_0_avalon_scaler_source_ready = video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module video_vga_controller_0_avalon_vga_sink_arbitrator (
                                                           // inputs:
                                                            clk,
                                                            reset_n,
                                                            video_dual_clock_buffer_0_avalon_dc_buffer_source_data,
                                                            video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket,
                                                            video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket,
                                                            video_dual_clock_buffer_0_avalon_dc_buffer_source_valid,
                                                            video_vga_controller_0_avalon_vga_sink_ready,

                                                           // outputs:
                                                            video_vga_controller_0_avalon_vga_sink_data,
                                                            video_vga_controller_0_avalon_vga_sink_endofpacket,
                                                            video_vga_controller_0_avalon_vga_sink_ready_from_sa,
                                                            video_vga_controller_0_avalon_vga_sink_reset,
                                                            video_vga_controller_0_avalon_vga_sink_startofpacket,
                                                            video_vga_controller_0_avalon_vga_sink_valid
                                                         )
;

  output  [ 29: 0] video_vga_controller_0_avalon_vga_sink_data;
  output           video_vga_controller_0_avalon_vga_sink_endofpacket;
  output           video_vga_controller_0_avalon_vga_sink_ready_from_sa;
  output           video_vga_controller_0_avalon_vga_sink_reset;
  output           video_vga_controller_0_avalon_vga_sink_startofpacket;
  output           video_vga_controller_0_avalon_vga_sink_valid;
  input            clk;
  input            reset_n;
  input   [ 29: 0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;
  input            video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;
  input            video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;
  input            video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;
  input            video_vga_controller_0_avalon_vga_sink_ready;

  wire    [ 29: 0] video_vga_controller_0_avalon_vga_sink_data;
  wire             video_vga_controller_0_avalon_vga_sink_endofpacket;
  wire             video_vga_controller_0_avalon_vga_sink_ready_from_sa;
  wire             video_vga_controller_0_avalon_vga_sink_reset;
  wire             video_vga_controller_0_avalon_vga_sink_startofpacket;
  wire             video_vga_controller_0_avalon_vga_sink_valid;
  //mux video_vga_controller_0_avalon_vga_sink_data, which is an e_mux
  assign video_vga_controller_0_avalon_vga_sink_data = video_dual_clock_buffer_0_avalon_dc_buffer_source_data;

  //mux video_vga_controller_0_avalon_vga_sink_endofpacket, which is an e_mux
  assign video_vga_controller_0_avalon_vga_sink_endofpacket = video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;

  //assign video_vga_controller_0_avalon_vga_sink_ready_from_sa = video_vga_controller_0_avalon_vga_sink_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign video_vga_controller_0_avalon_vga_sink_ready_from_sa = video_vga_controller_0_avalon_vga_sink_ready;

  //mux video_vga_controller_0_avalon_vga_sink_startofpacket, which is an e_mux
  assign video_vga_controller_0_avalon_vga_sink_startofpacket = video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;

  //mux video_vga_controller_0_avalon_vga_sink_valid, which is an e_mux
  assign video_vga_controller_0_avalon_vga_sink_valid = video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;

  //~video_vga_controller_0_avalon_vga_sink_reset assignment, which is an e_assign
  assign video_vga_controller_0_avalon_vga_sink_reset = ~reset_n;


endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_reset_clk_0_domain_synch_module (
                                                     // inputs:
                                                      clk,
                                                      data_in,
                                                      reset_n,

                                                     // outputs:
                                                      data_out
                                                   )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_reset_sys_clk_domain_synch_module (
                                                       // inputs:
                                                        clk,
                                                        data_in,
                                                        reset_n,

                                                       // outputs:
                                                        data_out
                                                     )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_reset_sdram_clk_domain_synch_module (
                                                         // inputs:
                                                          clk,
                                                          data_in,
                                                          reset_n,

                                                         // outputs:
                                                          data_out
                                                       )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system_reset_vga_clock_domain_synch_module (
                                                         // inputs:
                                                          clk,
                                                          data_in,
                                                          reset_n,

                                                         // outputs:
                                                          data_out
                                                       )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule


// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nios_system (
                     // 1) global signals:
                      clk_0,
                      reset_n,
                      sdram_clk,
                      sys_clk,
                      vga_clock,

                     // the_keys
                      in_port_to_the_keys,

                     // the_sdram_0
                      zs_addr_from_the_sdram_0,
                      zs_ba_from_the_sdram_0,
                      zs_cas_n_from_the_sdram_0,
                      zs_cke_from_the_sdram_0,
                      zs_cs_n_from_the_sdram_0,
                      zs_dq_to_and_from_the_sdram_0,
                      zs_dqm_from_the_sdram_0,
                      zs_ras_n_from_the_sdram_0,
                      zs_we_n_from_the_sdram_0,

                     // the_sram_0
                      SRAM_ADDR_from_the_sram_0,
                      SRAM_CE_N_from_the_sram_0,
                      SRAM_DQ_to_and_from_the_sram_0,
                      SRAM_LB_N_from_the_sram_0,
                      SRAM_OE_N_from_the_sram_0,
                      SRAM_UB_N_from_the_sram_0,
                      SRAM_WE_N_from_the_sram_0,

                     // the_video_vga_controller_0
                      VGA_BLANK_from_the_video_vga_controller_0,
                      VGA_B_from_the_video_vga_controller_0,
                      VGA_CLK_from_the_video_vga_controller_0,
                      VGA_G_from_the_video_vga_controller_0,
                      VGA_HS_from_the_video_vga_controller_0,
                      VGA_R_from_the_video_vga_controller_0,
                      VGA_SYNC_from_the_video_vga_controller_0,
                      VGA_VS_from_the_video_vga_controller_0
                   )
;

  output  [ 17: 0] SRAM_ADDR_from_the_sram_0;
  output           SRAM_CE_N_from_the_sram_0;
  inout   [ 15: 0] SRAM_DQ_to_and_from_the_sram_0;
  output           SRAM_LB_N_from_the_sram_0;
  output           SRAM_OE_N_from_the_sram_0;
  output           SRAM_UB_N_from_the_sram_0;
  output           SRAM_WE_N_from_the_sram_0;
  output           VGA_BLANK_from_the_video_vga_controller_0;
  output  [  9: 0] VGA_B_from_the_video_vga_controller_0;
  output           VGA_CLK_from_the_video_vga_controller_0;
  output  [  9: 0] VGA_G_from_the_video_vga_controller_0;
  output           VGA_HS_from_the_video_vga_controller_0;
  output  [  9: 0] VGA_R_from_the_video_vga_controller_0;
  output           VGA_SYNC_from_the_video_vga_controller_0;
  output           VGA_VS_from_the_video_vga_controller_0;
  output           sdram_clk;
  output           sys_clk;
  output           vga_clock;
  output  [ 11: 0] zs_addr_from_the_sdram_0;
  output  [  1: 0] zs_ba_from_the_sdram_0;
  output           zs_cas_n_from_the_sdram_0;
  output           zs_cke_from_the_sdram_0;
  output           zs_cs_n_from_the_sdram_0;
  inout   [ 15: 0] zs_dq_to_and_from_the_sdram_0;
  output  [  1: 0] zs_dqm_from_the_sdram_0;
  output           zs_ras_n_from_the_sdram_0;
  output           zs_we_n_from_the_sdram_0;
  input            clk_0;
  input   [  2: 0] in_port_to_the_keys;
  input            reset_n;

  wire    [ 17: 0] SRAM_ADDR_from_the_sram_0;
  wire             SRAM_CE_N_from_the_sram_0;
  wire    [ 15: 0] SRAM_DQ_to_and_from_the_sram_0;
  wire             SRAM_LB_N_from_the_sram_0;
  wire             SRAM_OE_N_from_the_sram_0;
  wire             SRAM_UB_N_from_the_sram_0;
  wire             SRAM_WE_N_from_the_sram_0;
  wire             VGA_BLANK_from_the_video_vga_controller_0;
  wire    [  9: 0] VGA_B_from_the_video_vga_controller_0;
  wire             VGA_CLK_from_the_video_vga_controller_0;
  wire    [  9: 0] VGA_G_from_the_video_vga_controller_0;
  wire             VGA_HS_from_the_video_vga_controller_0;
  wire    [  9: 0] VGA_R_from_the_video_vga_controller_0;
  wire             VGA_SYNC_from_the_video_vga_controller_0;
  wire             VGA_VS_from_the_video_vga_controller_0;
  wire             clk_0_reset_n;
  wire             clocks_0_avalon_clocks_slave_address;
  wire    [  7: 0] clocks_0_avalon_clocks_slave_readdata;
  wire    [  7: 0] clocks_0_avalon_clocks_slave_readdata_from_sa;
  wire             cpu_0_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  wire    [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  wire    [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_datab;
  wire             cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done;
  wire             cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  wire    [  1: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_n;
  wire             cpu_0_altera_nios_custom_instr_floating_point_inst_s1_reset;
  wire    [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result;
  wire    [ 31: 0] cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  wire             cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select;
  wire             cpu_0_altera_nios_custom_instr_floating_point_inst_s1_start;
  wire    [  4: 0] cpu_0_custom_instruction_master_multi_a;
  wire    [  4: 0] cpu_0_custom_instruction_master_multi_b;
  wire    [  4: 0] cpu_0_custom_instruction_master_multi_c;
  wire             cpu_0_custom_instruction_master_multi_clk;
  wire             cpu_0_custom_instruction_master_multi_clk_en;
  wire    [ 31: 0] cpu_0_custom_instruction_master_multi_dataa;
  wire    [ 31: 0] cpu_0_custom_instruction_master_multi_datab;
  wire             cpu_0_custom_instruction_master_multi_done;
  wire             cpu_0_custom_instruction_master_multi_estatus;
  wire    [ 31: 0] cpu_0_custom_instruction_master_multi_ipending;
  wire    [  7: 0] cpu_0_custom_instruction_master_multi_n;
  wire             cpu_0_custom_instruction_master_multi_readra;
  wire             cpu_0_custom_instruction_master_multi_readrb;
  wire             cpu_0_custom_instruction_master_multi_reset;
  wire    [ 31: 0] cpu_0_custom_instruction_master_multi_result;
  wire             cpu_0_custom_instruction_master_multi_start;
  wire             cpu_0_custom_instruction_master_multi_status;
  wire             cpu_0_custom_instruction_master_multi_writerc;
  wire             cpu_0_custom_instruction_master_reset_n;
  wire             cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1;
  wire    [ 24: 0] cpu_0_data_master_address;
  wire    [ 24: 0] cpu_0_data_master_address_to_slave;
  wire    [  3: 0] cpu_0_data_master_byteenable;
  wire    [  1: 0] cpu_0_data_master_byteenable_nios_system_clock_3_in;
  wire             cpu_0_data_master_byteenable_nios_system_clock_9_in;
  wire    [  1: 0] cpu_0_data_master_byteenable_sram_0_avalon_sram_slave;
  wire    [  1: 0] cpu_0_data_master_dbs_address;
  wire    [ 15: 0] cpu_0_data_master_dbs_write_16;
  wire    [  7: 0] cpu_0_data_master_dbs_write_8;
  wire             cpu_0_data_master_debugaccess;
  wire             cpu_0_data_master_granted_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_granted_keys_s1;
  wire             cpu_0_data_master_granted_mailbox_0_s1;
  wire             cpu_0_data_master_granted_mailbox_1_s1;
  wire             cpu_0_data_master_granted_mailbox_2_s1;
  wire             cpu_0_data_master_granted_mailbox_3_s1;
  wire             cpu_0_data_master_granted_nios_system_clock_3_in;
  wire             cpu_0_data_master_granted_nios_system_clock_9_in;
  wire             cpu_0_data_master_granted_onchip_memory2_0_s1;
  wire             cpu_0_data_master_granted_onchip_memory2_1_s1;
  wire             cpu_0_data_master_granted_onchip_memory2_2_s1;
  wire             cpu_0_data_master_granted_onchip_memory2_3_s1;
  wire             cpu_0_data_master_granted_performance_counter_0_control_slave;
  wire             cpu_0_data_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_0_data_master_granted_sysid_control_slave;
  wire             cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  wire    [ 31: 0] cpu_0_data_master_irq;
  wire             cpu_0_data_master_latency_counter;
  wire             cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_qualified_request_keys_s1;
  wire             cpu_0_data_master_qualified_request_mailbox_0_s1;
  wire             cpu_0_data_master_qualified_request_mailbox_1_s1;
  wire             cpu_0_data_master_qualified_request_mailbox_2_s1;
  wire             cpu_0_data_master_qualified_request_mailbox_3_s1;
  wire             cpu_0_data_master_qualified_request_nios_system_clock_3_in;
  wire             cpu_0_data_master_qualified_request_nios_system_clock_9_in;
  wire             cpu_0_data_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_0_data_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_0_data_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_0_data_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_0_data_master_qualified_request_performance_counter_0_control_slave;
  wire             cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_0_data_master_qualified_request_sysid_control_slave;
  wire             cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_0_data_master_read;
  wire             cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_read_data_valid_keys_s1;
  wire             cpu_0_data_master_read_data_valid_mailbox_0_s1;
  wire             cpu_0_data_master_read_data_valid_mailbox_1_s1;
  wire             cpu_0_data_master_read_data_valid_mailbox_2_s1;
  wire             cpu_0_data_master_read_data_valid_mailbox_3_s1;
  wire             cpu_0_data_master_read_data_valid_nios_system_clock_3_in;
  wire             cpu_0_data_master_read_data_valid_nios_system_clock_9_in;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_0_s1;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_1_s1;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_2_s1;
  wire             cpu_0_data_master_read_data_valid_onchip_memory2_3_s1;
  wire             cpu_0_data_master_read_data_valid_performance_counter_0_control_slave;
  wire             cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             cpu_0_data_master_read_data_valid_sysid_control_slave;
  wire             cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  wire    [ 31: 0] cpu_0_data_master_readdata;
  wire             cpu_0_data_master_readdatavalid;
  wire             cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_requests_keys_s1;
  wire             cpu_0_data_master_requests_mailbox_0_s1;
  wire             cpu_0_data_master_requests_mailbox_1_s1;
  wire             cpu_0_data_master_requests_mailbox_2_s1;
  wire             cpu_0_data_master_requests_mailbox_3_s1;
  wire             cpu_0_data_master_requests_nios_system_clock_3_in;
  wire             cpu_0_data_master_requests_nios_system_clock_9_in;
  wire             cpu_0_data_master_requests_onchip_memory2_0_s1;
  wire             cpu_0_data_master_requests_onchip_memory2_1_s1;
  wire             cpu_0_data_master_requests_onchip_memory2_2_s1;
  wire             cpu_0_data_master_requests_onchip_memory2_3_s1;
  wire             cpu_0_data_master_requests_performance_counter_0_control_slave;
  wire             cpu_0_data_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_0_data_master_requests_sysid_control_slave;
  wire             cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_0_data_master_waitrequest;
  wire             cpu_0_data_master_write;
  wire    [ 31: 0] cpu_0_data_master_writedata;
  wire    [ 24: 0] cpu_0_instruction_master_address;
  wire    [ 24: 0] cpu_0_instruction_master_address_to_slave;
  wire    [  1: 0] cpu_0_instruction_master_dbs_address;
  wire             cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_granted_nios_system_clock_2_in;
  wire             cpu_0_instruction_master_granted_onchip_memory2_0_s1;
  wire             cpu_0_instruction_master_granted_onchip_memory2_1_s1;
  wire             cpu_0_instruction_master_granted_onchip_memory2_2_s1;
  wire             cpu_0_instruction_master_granted_onchip_memory2_3_s1;
  wire             cpu_0_instruction_master_latency_counter;
  wire             cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_qualified_request_nios_system_clock_2_in;
  wire             cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_0_instruction_master_read;
  wire             cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1;
  wire             cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1;
  wire    [ 31: 0] cpu_0_instruction_master_readdata;
  wire             cpu_0_instruction_master_readdatavalid;
  wire             cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_requests_nios_system_clock_2_in;
  wire             cpu_0_instruction_master_requests_onchip_memory2_0_s1;
  wire             cpu_0_instruction_master_requests_onchip_memory2_1_s1;
  wire             cpu_0_instruction_master_requests_onchip_memory2_2_s1;
  wire             cpu_0_instruction_master_requests_onchip_memory2_3_s1;
  wire             cpu_0_instruction_master_waitrequest;
  wire    [  8: 0] cpu_0_jtag_debug_module_address;
  wire             cpu_0_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_0_jtag_debug_module_byteenable;
  wire             cpu_0_jtag_debug_module_chipselect;
  wire             cpu_0_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_0_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_0_jtag_debug_module_readdata_from_sa;
  wire             cpu_0_jtag_debug_module_resetrequest;
  wire             cpu_0_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_0_jtag_debug_module_write;
  wire    [ 31: 0] cpu_0_jtag_debug_module_writedata;
  wire             cpu_1_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  wire    [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  wire    [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_datab;
  wire             cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done;
  wire             cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  wire    [  1: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_n;
  wire             cpu_1_altera_nios_custom_instr_floating_point_inst_s1_reset;
  wire    [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result;
  wire    [ 31: 0] cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  wire             cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select;
  wire             cpu_1_altera_nios_custom_instr_floating_point_inst_s1_start;
  wire    [  4: 0] cpu_1_custom_instruction_master_multi_a;
  wire    [  4: 0] cpu_1_custom_instruction_master_multi_b;
  wire    [  4: 0] cpu_1_custom_instruction_master_multi_c;
  wire             cpu_1_custom_instruction_master_multi_clk;
  wire             cpu_1_custom_instruction_master_multi_clk_en;
  wire    [ 31: 0] cpu_1_custom_instruction_master_multi_dataa;
  wire    [ 31: 0] cpu_1_custom_instruction_master_multi_datab;
  wire             cpu_1_custom_instruction_master_multi_done;
  wire             cpu_1_custom_instruction_master_multi_estatus;
  wire    [ 31: 0] cpu_1_custom_instruction_master_multi_ipending;
  wire    [  7: 0] cpu_1_custom_instruction_master_multi_n;
  wire             cpu_1_custom_instruction_master_multi_readra;
  wire             cpu_1_custom_instruction_master_multi_readrb;
  wire             cpu_1_custom_instruction_master_multi_reset;
  wire    [ 31: 0] cpu_1_custom_instruction_master_multi_result;
  wire             cpu_1_custom_instruction_master_multi_start;
  wire             cpu_1_custom_instruction_master_multi_status;
  wire             cpu_1_custom_instruction_master_multi_writerc;
  wire             cpu_1_custom_instruction_master_reset_n;
  wire             cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1;
  wire    [ 24: 0] cpu_1_data_master_address;
  wire    [ 24: 0] cpu_1_data_master_address_to_slave;
  wire    [  3: 0] cpu_1_data_master_byteenable;
  wire    [  1: 0] cpu_1_data_master_byteenable_nios_system_clock_1_in;
  wire             cpu_1_data_master_byteenable_nios_system_clock_8_in;
  wire    [  1: 0] cpu_1_data_master_byteenable_sram_0_avalon_sram_slave;
  wire    [  1: 0] cpu_1_data_master_dbs_address;
  wire    [ 15: 0] cpu_1_data_master_dbs_write_16;
  wire    [  7: 0] cpu_1_data_master_dbs_write_8;
  wire             cpu_1_data_master_debugaccess;
  wire             cpu_1_data_master_granted_cpu_1_jtag_debug_module;
  wire             cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave;
  wire             cpu_1_data_master_granted_keys_s1;
  wire             cpu_1_data_master_granted_mailbox_0_s1;
  wire             cpu_1_data_master_granted_mailbox_1_s1;
  wire             cpu_1_data_master_granted_mailbox_2_s1;
  wire             cpu_1_data_master_granted_mailbox_3_s1;
  wire             cpu_1_data_master_granted_nios_system_clock_1_in;
  wire             cpu_1_data_master_granted_nios_system_clock_8_in;
  wire             cpu_1_data_master_granted_onchip_memory2_0_s1;
  wire             cpu_1_data_master_granted_onchip_memory2_1_s1;
  wire             cpu_1_data_master_granted_onchip_memory2_2_s1;
  wire             cpu_1_data_master_granted_onchip_memory2_3_s1;
  wire             cpu_1_data_master_granted_performance_counter_0_control_slave;
  wire             cpu_1_data_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_1_data_master_granted_sysid_control_slave;
  wire             cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  wire    [ 31: 0] cpu_1_data_master_irq;
  wire             cpu_1_data_master_latency_counter;
  wire             cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module;
  wire             cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave;
  wire             cpu_1_data_master_qualified_request_keys_s1;
  wire             cpu_1_data_master_qualified_request_mailbox_0_s1;
  wire             cpu_1_data_master_qualified_request_mailbox_1_s1;
  wire             cpu_1_data_master_qualified_request_mailbox_2_s1;
  wire             cpu_1_data_master_qualified_request_mailbox_3_s1;
  wire             cpu_1_data_master_qualified_request_nios_system_clock_1_in;
  wire             cpu_1_data_master_qualified_request_nios_system_clock_8_in;
  wire             cpu_1_data_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_1_data_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_1_data_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_1_data_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_1_data_master_qualified_request_performance_counter_0_control_slave;
  wire             cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_1_data_master_qualified_request_sysid_control_slave;
  wire             cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_1_data_master_read;
  wire             cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module;
  wire             cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave;
  wire             cpu_1_data_master_read_data_valid_keys_s1;
  wire             cpu_1_data_master_read_data_valid_mailbox_0_s1;
  wire             cpu_1_data_master_read_data_valid_mailbox_1_s1;
  wire             cpu_1_data_master_read_data_valid_mailbox_2_s1;
  wire             cpu_1_data_master_read_data_valid_mailbox_3_s1;
  wire             cpu_1_data_master_read_data_valid_nios_system_clock_1_in;
  wire             cpu_1_data_master_read_data_valid_nios_system_clock_8_in;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_0_s1;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_1_s1;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_2_s1;
  wire             cpu_1_data_master_read_data_valid_onchip_memory2_3_s1;
  wire             cpu_1_data_master_read_data_valid_performance_counter_0_control_slave;
  wire             cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             cpu_1_data_master_read_data_valid_sysid_control_slave;
  wire             cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  wire    [ 31: 0] cpu_1_data_master_readdata;
  wire             cpu_1_data_master_readdatavalid;
  wire             cpu_1_data_master_requests_cpu_1_jtag_debug_module;
  wire             cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave;
  wire             cpu_1_data_master_requests_keys_s1;
  wire             cpu_1_data_master_requests_mailbox_0_s1;
  wire             cpu_1_data_master_requests_mailbox_1_s1;
  wire             cpu_1_data_master_requests_mailbox_2_s1;
  wire             cpu_1_data_master_requests_mailbox_3_s1;
  wire             cpu_1_data_master_requests_nios_system_clock_1_in;
  wire             cpu_1_data_master_requests_nios_system_clock_8_in;
  wire             cpu_1_data_master_requests_onchip_memory2_0_s1;
  wire             cpu_1_data_master_requests_onchip_memory2_1_s1;
  wire             cpu_1_data_master_requests_onchip_memory2_2_s1;
  wire             cpu_1_data_master_requests_onchip_memory2_3_s1;
  wire             cpu_1_data_master_requests_performance_counter_0_control_slave;
  wire             cpu_1_data_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_1_data_master_requests_sysid_control_slave;
  wire             cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_1_data_master_waitrequest;
  wire             cpu_1_data_master_write;
  wire    [ 31: 0] cpu_1_data_master_writedata;
  wire    [ 24: 0] cpu_1_instruction_master_address;
  wire    [ 24: 0] cpu_1_instruction_master_address_to_slave;
  wire    [  1: 0] cpu_1_instruction_master_dbs_address;
  wire             cpu_1_instruction_master_granted_cpu_1_jtag_debug_module;
  wire             cpu_1_instruction_master_granted_nios_system_clock_0_in;
  wire             cpu_1_instruction_master_granted_onchip_memory2_0_s1;
  wire             cpu_1_instruction_master_granted_onchip_memory2_1_s1;
  wire             cpu_1_instruction_master_granted_onchip_memory2_2_s1;
  wire             cpu_1_instruction_master_granted_onchip_memory2_3_s1;
  wire             cpu_1_instruction_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_1_instruction_master_latency_counter;
  wire             cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module;
  wire             cpu_1_instruction_master_qualified_request_nios_system_clock_0_in;
  wire             cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_1_instruction_master_read;
  wire             cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module;
  wire             cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1;
  wire             cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1;
  wire             cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire    [ 31: 0] cpu_1_instruction_master_readdata;
  wire             cpu_1_instruction_master_readdatavalid;
  wire             cpu_1_instruction_master_requests_cpu_1_jtag_debug_module;
  wire             cpu_1_instruction_master_requests_nios_system_clock_0_in;
  wire             cpu_1_instruction_master_requests_onchip_memory2_0_s1;
  wire             cpu_1_instruction_master_requests_onchip_memory2_1_s1;
  wire             cpu_1_instruction_master_requests_onchip_memory2_2_s1;
  wire             cpu_1_instruction_master_requests_onchip_memory2_3_s1;
  wire             cpu_1_instruction_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_1_instruction_master_waitrequest;
  wire    [  8: 0] cpu_1_jtag_debug_module_address;
  wire             cpu_1_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_1_jtag_debug_module_byteenable;
  wire             cpu_1_jtag_debug_module_chipselect;
  wire             cpu_1_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_1_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_1_jtag_debug_module_readdata_from_sa;
  wire             cpu_1_jtag_debug_module_resetrequest;
  wire             cpu_1_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_1_jtag_debug_module_write;
  wire    [ 31: 0] cpu_1_jtag_debug_module_writedata;
  wire             cpu_2_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  wire    [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  wire    [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_datab;
  wire             cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done;
  wire             cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  wire    [  1: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_n;
  wire             cpu_2_altera_nios_custom_instr_floating_point_inst_s1_reset;
  wire    [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result;
  wire    [ 31: 0] cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  wire             cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select;
  wire             cpu_2_altera_nios_custom_instr_floating_point_inst_s1_start;
  wire    [  4: 0] cpu_2_custom_instruction_master_multi_a;
  wire    [  4: 0] cpu_2_custom_instruction_master_multi_b;
  wire    [  4: 0] cpu_2_custom_instruction_master_multi_c;
  wire             cpu_2_custom_instruction_master_multi_clk;
  wire             cpu_2_custom_instruction_master_multi_clk_en;
  wire    [ 31: 0] cpu_2_custom_instruction_master_multi_dataa;
  wire    [ 31: 0] cpu_2_custom_instruction_master_multi_datab;
  wire             cpu_2_custom_instruction_master_multi_done;
  wire             cpu_2_custom_instruction_master_multi_estatus;
  wire    [ 31: 0] cpu_2_custom_instruction_master_multi_ipending;
  wire    [  7: 0] cpu_2_custom_instruction_master_multi_n;
  wire             cpu_2_custom_instruction_master_multi_readra;
  wire             cpu_2_custom_instruction_master_multi_readrb;
  wire             cpu_2_custom_instruction_master_multi_reset;
  wire    [ 31: 0] cpu_2_custom_instruction_master_multi_result;
  wire             cpu_2_custom_instruction_master_multi_start;
  wire             cpu_2_custom_instruction_master_multi_status;
  wire             cpu_2_custom_instruction_master_multi_writerc;
  wire             cpu_2_custom_instruction_master_reset_n;
  wire             cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1;
  wire    [ 24: 0] cpu_2_data_master_address;
  wire    [ 24: 0] cpu_2_data_master_address_to_slave;
  wire    [  3: 0] cpu_2_data_master_byteenable;
  wire             cpu_2_data_master_byteenable_nios_system_clock_10_in;
  wire    [  1: 0] cpu_2_data_master_byteenable_nios_system_clock_5_in;
  wire    [  1: 0] cpu_2_data_master_byteenable_sram_0_avalon_sram_slave;
  wire    [  1: 0] cpu_2_data_master_dbs_address;
  wire    [ 15: 0] cpu_2_data_master_dbs_write_16;
  wire    [  7: 0] cpu_2_data_master_dbs_write_8;
  wire             cpu_2_data_master_debugaccess;
  wire             cpu_2_data_master_granted_cpu_2_jtag_debug_module;
  wire             cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave;
  wire             cpu_2_data_master_granted_keys_s1;
  wire             cpu_2_data_master_granted_mailbox_0_s1;
  wire             cpu_2_data_master_granted_mailbox_1_s1;
  wire             cpu_2_data_master_granted_mailbox_2_s1;
  wire             cpu_2_data_master_granted_mailbox_3_s1;
  wire             cpu_2_data_master_granted_nios_system_clock_10_in;
  wire             cpu_2_data_master_granted_nios_system_clock_5_in;
  wire             cpu_2_data_master_granted_onchip_memory2_0_s1;
  wire             cpu_2_data_master_granted_onchip_memory2_1_s1;
  wire             cpu_2_data_master_granted_onchip_memory2_2_s1;
  wire             cpu_2_data_master_granted_onchip_memory2_3_s1;
  wire             cpu_2_data_master_granted_performance_counter_0_control_slave;
  wire             cpu_2_data_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_2_data_master_granted_sysid_control_slave;
  wire             cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  wire    [ 31: 0] cpu_2_data_master_irq;
  wire             cpu_2_data_master_latency_counter;
  wire             cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module;
  wire             cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave;
  wire             cpu_2_data_master_qualified_request_keys_s1;
  wire             cpu_2_data_master_qualified_request_mailbox_0_s1;
  wire             cpu_2_data_master_qualified_request_mailbox_1_s1;
  wire             cpu_2_data_master_qualified_request_mailbox_2_s1;
  wire             cpu_2_data_master_qualified_request_mailbox_3_s1;
  wire             cpu_2_data_master_qualified_request_nios_system_clock_10_in;
  wire             cpu_2_data_master_qualified_request_nios_system_clock_5_in;
  wire             cpu_2_data_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_2_data_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_2_data_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_2_data_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_2_data_master_qualified_request_performance_counter_0_control_slave;
  wire             cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_2_data_master_qualified_request_sysid_control_slave;
  wire             cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_2_data_master_read;
  wire             cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module;
  wire             cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave;
  wire             cpu_2_data_master_read_data_valid_keys_s1;
  wire             cpu_2_data_master_read_data_valid_mailbox_0_s1;
  wire             cpu_2_data_master_read_data_valid_mailbox_1_s1;
  wire             cpu_2_data_master_read_data_valid_mailbox_2_s1;
  wire             cpu_2_data_master_read_data_valid_mailbox_3_s1;
  wire             cpu_2_data_master_read_data_valid_nios_system_clock_10_in;
  wire             cpu_2_data_master_read_data_valid_nios_system_clock_5_in;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_0_s1;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_1_s1;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_2_s1;
  wire             cpu_2_data_master_read_data_valid_onchip_memory2_3_s1;
  wire             cpu_2_data_master_read_data_valid_performance_counter_0_control_slave;
  wire             cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             cpu_2_data_master_read_data_valid_sysid_control_slave;
  wire             cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  wire    [ 31: 0] cpu_2_data_master_readdata;
  wire             cpu_2_data_master_readdatavalid;
  wire             cpu_2_data_master_requests_cpu_2_jtag_debug_module;
  wire             cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave;
  wire             cpu_2_data_master_requests_keys_s1;
  wire             cpu_2_data_master_requests_mailbox_0_s1;
  wire             cpu_2_data_master_requests_mailbox_1_s1;
  wire             cpu_2_data_master_requests_mailbox_2_s1;
  wire             cpu_2_data_master_requests_mailbox_3_s1;
  wire             cpu_2_data_master_requests_nios_system_clock_10_in;
  wire             cpu_2_data_master_requests_nios_system_clock_5_in;
  wire             cpu_2_data_master_requests_onchip_memory2_0_s1;
  wire             cpu_2_data_master_requests_onchip_memory2_1_s1;
  wire             cpu_2_data_master_requests_onchip_memory2_2_s1;
  wire             cpu_2_data_master_requests_onchip_memory2_3_s1;
  wire             cpu_2_data_master_requests_performance_counter_0_control_slave;
  wire             cpu_2_data_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_2_data_master_requests_sysid_control_slave;
  wire             cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_2_data_master_waitrequest;
  wire             cpu_2_data_master_write;
  wire    [ 31: 0] cpu_2_data_master_writedata;
  wire    [ 24: 0] cpu_2_instruction_master_address;
  wire    [ 24: 0] cpu_2_instruction_master_address_to_slave;
  wire    [  1: 0] cpu_2_instruction_master_dbs_address;
  wire             cpu_2_instruction_master_granted_cpu_2_jtag_debug_module;
  wire             cpu_2_instruction_master_granted_nios_system_clock_4_in;
  wire             cpu_2_instruction_master_granted_onchip_memory2_0_s1;
  wire             cpu_2_instruction_master_granted_onchip_memory2_1_s1;
  wire             cpu_2_instruction_master_granted_onchip_memory2_2_s1;
  wire             cpu_2_instruction_master_granted_onchip_memory2_3_s1;
  wire             cpu_2_instruction_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_2_instruction_master_latency_counter;
  wire             cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module;
  wire             cpu_2_instruction_master_qualified_request_nios_system_clock_4_in;
  wire             cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_2_instruction_master_read;
  wire             cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module;
  wire             cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1;
  wire             cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1;
  wire             cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire    [ 31: 0] cpu_2_instruction_master_readdata;
  wire             cpu_2_instruction_master_readdatavalid;
  wire             cpu_2_instruction_master_requests_cpu_2_jtag_debug_module;
  wire             cpu_2_instruction_master_requests_nios_system_clock_4_in;
  wire             cpu_2_instruction_master_requests_onchip_memory2_0_s1;
  wire             cpu_2_instruction_master_requests_onchip_memory2_1_s1;
  wire             cpu_2_instruction_master_requests_onchip_memory2_2_s1;
  wire             cpu_2_instruction_master_requests_onchip_memory2_3_s1;
  wire             cpu_2_instruction_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_2_instruction_master_waitrequest;
  wire    [  8: 0] cpu_2_jtag_debug_module_address;
  wire             cpu_2_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_2_jtag_debug_module_byteenable;
  wire             cpu_2_jtag_debug_module_chipselect;
  wire             cpu_2_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_2_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_2_jtag_debug_module_readdata_from_sa;
  wire             cpu_2_jtag_debug_module_resetrequest;
  wire             cpu_2_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_2_jtag_debug_module_write;
  wire    [ 31: 0] cpu_2_jtag_debug_module_writedata;
  wire             cpu_3_altera_nios_custom_instr_floating_point_inst_s1_clk_en;
  wire    [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_dataa;
  wire    [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_datab;
  wire             cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done;
  wire             cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa;
  wire    [  1: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_n;
  wire             cpu_3_altera_nios_custom_instr_floating_point_inst_s1_reset;
  wire    [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result;
  wire    [ 31: 0] cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa;
  wire             cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select;
  wire             cpu_3_altera_nios_custom_instr_floating_point_inst_s1_start;
  wire    [  4: 0] cpu_3_custom_instruction_master_multi_a;
  wire    [  4: 0] cpu_3_custom_instruction_master_multi_b;
  wire    [  4: 0] cpu_3_custom_instruction_master_multi_c;
  wire             cpu_3_custom_instruction_master_multi_clk;
  wire             cpu_3_custom_instruction_master_multi_clk_en;
  wire    [ 31: 0] cpu_3_custom_instruction_master_multi_dataa;
  wire    [ 31: 0] cpu_3_custom_instruction_master_multi_datab;
  wire             cpu_3_custom_instruction_master_multi_done;
  wire             cpu_3_custom_instruction_master_multi_estatus;
  wire    [ 31: 0] cpu_3_custom_instruction_master_multi_ipending;
  wire    [  7: 0] cpu_3_custom_instruction_master_multi_n;
  wire             cpu_3_custom_instruction_master_multi_readra;
  wire             cpu_3_custom_instruction_master_multi_readrb;
  wire             cpu_3_custom_instruction_master_multi_reset;
  wire    [ 31: 0] cpu_3_custom_instruction_master_multi_result;
  wire             cpu_3_custom_instruction_master_multi_start;
  wire             cpu_3_custom_instruction_master_multi_status;
  wire             cpu_3_custom_instruction_master_multi_writerc;
  wire             cpu_3_custom_instruction_master_reset_n;
  wire             cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1;
  wire    [ 24: 0] cpu_3_data_master_address;
  wire    [ 24: 0] cpu_3_data_master_address_to_slave;
  wire    [  3: 0] cpu_3_data_master_byteenable;
  wire             cpu_3_data_master_byteenable_nios_system_clock_11_in;
  wire    [  1: 0] cpu_3_data_master_byteenable_nios_system_clock_7_in;
  wire    [  1: 0] cpu_3_data_master_byteenable_sram_0_avalon_sram_slave;
  wire    [  1: 0] cpu_3_data_master_dbs_address;
  wire    [ 15: 0] cpu_3_data_master_dbs_write_16;
  wire    [  7: 0] cpu_3_data_master_dbs_write_8;
  wire             cpu_3_data_master_debugaccess;
  wire             cpu_3_data_master_granted_cpu_3_jtag_debug_module;
  wire             cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave;
  wire             cpu_3_data_master_granted_keys_s1;
  wire             cpu_3_data_master_granted_mailbox_0_s1;
  wire             cpu_3_data_master_granted_mailbox_1_s1;
  wire             cpu_3_data_master_granted_mailbox_2_s1;
  wire             cpu_3_data_master_granted_mailbox_3_s1;
  wire             cpu_3_data_master_granted_nios_system_clock_11_in;
  wire             cpu_3_data_master_granted_nios_system_clock_7_in;
  wire             cpu_3_data_master_granted_onchip_memory2_0_s1;
  wire             cpu_3_data_master_granted_onchip_memory2_1_s1;
  wire             cpu_3_data_master_granted_onchip_memory2_2_s1;
  wire             cpu_3_data_master_granted_onchip_memory2_3_s1;
  wire             cpu_3_data_master_granted_performance_counter_0_control_slave;
  wire             cpu_3_data_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_3_data_master_granted_sysid_control_slave;
  wire             cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave;
  wire    [ 31: 0] cpu_3_data_master_irq;
  wire             cpu_3_data_master_latency_counter;
  wire             cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module;
  wire             cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave;
  wire             cpu_3_data_master_qualified_request_keys_s1;
  wire             cpu_3_data_master_qualified_request_mailbox_0_s1;
  wire             cpu_3_data_master_qualified_request_mailbox_1_s1;
  wire             cpu_3_data_master_qualified_request_mailbox_2_s1;
  wire             cpu_3_data_master_qualified_request_mailbox_3_s1;
  wire             cpu_3_data_master_qualified_request_nios_system_clock_11_in;
  wire             cpu_3_data_master_qualified_request_nios_system_clock_7_in;
  wire             cpu_3_data_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_3_data_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_3_data_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_3_data_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_3_data_master_qualified_request_performance_counter_0_control_slave;
  wire             cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_3_data_master_qualified_request_sysid_control_slave;
  wire             cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_3_data_master_read;
  wire             cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module;
  wire             cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave;
  wire             cpu_3_data_master_read_data_valid_keys_s1;
  wire             cpu_3_data_master_read_data_valid_mailbox_0_s1;
  wire             cpu_3_data_master_read_data_valid_mailbox_1_s1;
  wire             cpu_3_data_master_read_data_valid_mailbox_2_s1;
  wire             cpu_3_data_master_read_data_valid_mailbox_3_s1;
  wire             cpu_3_data_master_read_data_valid_nios_system_clock_11_in;
  wire             cpu_3_data_master_read_data_valid_nios_system_clock_7_in;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_0_s1;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_1_s1;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_2_s1;
  wire             cpu_3_data_master_read_data_valid_onchip_memory2_3_s1;
  wire             cpu_3_data_master_read_data_valid_performance_counter_0_control_slave;
  wire             cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire             cpu_3_data_master_read_data_valid_sysid_control_slave;
  wire             cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave;
  wire    [ 31: 0] cpu_3_data_master_readdata;
  wire             cpu_3_data_master_readdatavalid;
  wire             cpu_3_data_master_requests_cpu_3_jtag_debug_module;
  wire             cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave;
  wire             cpu_3_data_master_requests_keys_s1;
  wire             cpu_3_data_master_requests_mailbox_0_s1;
  wire             cpu_3_data_master_requests_mailbox_1_s1;
  wire             cpu_3_data_master_requests_mailbox_2_s1;
  wire             cpu_3_data_master_requests_mailbox_3_s1;
  wire             cpu_3_data_master_requests_nios_system_clock_11_in;
  wire             cpu_3_data_master_requests_nios_system_clock_7_in;
  wire             cpu_3_data_master_requests_onchip_memory2_0_s1;
  wire             cpu_3_data_master_requests_onchip_memory2_1_s1;
  wire             cpu_3_data_master_requests_onchip_memory2_2_s1;
  wire             cpu_3_data_master_requests_onchip_memory2_3_s1;
  wire             cpu_3_data_master_requests_performance_counter_0_control_slave;
  wire             cpu_3_data_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_3_data_master_requests_sysid_control_slave;
  wire             cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave;
  wire             cpu_3_data_master_waitrequest;
  wire             cpu_3_data_master_write;
  wire    [ 31: 0] cpu_3_data_master_writedata;
  wire    [ 24: 0] cpu_3_instruction_master_address;
  wire    [ 24: 0] cpu_3_instruction_master_address_to_slave;
  wire    [  1: 0] cpu_3_instruction_master_dbs_address;
  wire             cpu_3_instruction_master_granted_cpu_3_jtag_debug_module;
  wire             cpu_3_instruction_master_granted_nios_system_clock_6_in;
  wire             cpu_3_instruction_master_granted_onchip_memory2_0_s1;
  wire             cpu_3_instruction_master_granted_onchip_memory2_1_s1;
  wire             cpu_3_instruction_master_granted_onchip_memory2_2_s1;
  wire             cpu_3_instruction_master_granted_onchip_memory2_3_s1;
  wire             cpu_3_instruction_master_granted_sram_0_avalon_sram_slave;
  wire             cpu_3_instruction_master_latency_counter;
  wire             cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module;
  wire             cpu_3_instruction_master_qualified_request_nios_system_clock_6_in;
  wire             cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1;
  wire             cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1;
  wire             cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1;
  wire             cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1;
  wire             cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave;
  wire             cpu_3_instruction_master_read;
  wire             cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module;
  wire             cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1;
  wire             cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1;
  wire             cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire    [ 31: 0] cpu_3_instruction_master_readdata;
  wire             cpu_3_instruction_master_readdatavalid;
  wire             cpu_3_instruction_master_requests_cpu_3_jtag_debug_module;
  wire             cpu_3_instruction_master_requests_nios_system_clock_6_in;
  wire             cpu_3_instruction_master_requests_onchip_memory2_0_s1;
  wire             cpu_3_instruction_master_requests_onchip_memory2_1_s1;
  wire             cpu_3_instruction_master_requests_onchip_memory2_2_s1;
  wire             cpu_3_instruction_master_requests_onchip_memory2_3_s1;
  wire             cpu_3_instruction_master_requests_sram_0_avalon_sram_slave;
  wire             cpu_3_instruction_master_waitrequest;
  wire    [  8: 0] cpu_3_jtag_debug_module_address;
  wire             cpu_3_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_3_jtag_debug_module_byteenable;
  wire             cpu_3_jtag_debug_module_chipselect;
  wire             cpu_3_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_3_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_3_jtag_debug_module_readdata_from_sa;
  wire             cpu_3_jtag_debug_module_resetrequest;
  wire             cpu_3_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_3_jtag_debug_module_write;
  wire    [ 31: 0] cpu_3_jtag_debug_module_writedata;
  wire             d1_clocks_0_avalon_clocks_slave_end_xfer;
  wire             d1_cpu_0_jtag_debug_module_end_xfer;
  wire             d1_cpu_1_jtag_debug_module_end_xfer;
  wire             d1_cpu_2_jtag_debug_module_end_xfer;
  wire             d1_cpu_3_jtag_debug_module_end_xfer;
  wire             d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  wire             d1_jtag_uart_1_avalon_jtag_slave_end_xfer;
  wire             d1_jtag_uart_2_avalon_jtag_slave_end_xfer;
  wire             d1_jtag_uart_3_avalon_jtag_slave_end_xfer;
  wire             d1_keys_s1_end_xfer;
  wire             d1_mailbox_0_s1_end_xfer;
  wire             d1_mailbox_1_s1_end_xfer;
  wire             d1_mailbox_2_s1_end_xfer;
  wire             d1_mailbox_3_s1_end_xfer;
  wire             d1_nios_system_clock_0_in_end_xfer;
  wire             d1_nios_system_clock_10_in_end_xfer;
  wire             d1_nios_system_clock_11_in_end_xfer;
  wire             d1_nios_system_clock_1_in_end_xfer;
  wire             d1_nios_system_clock_2_in_end_xfer;
  wire             d1_nios_system_clock_3_in_end_xfer;
  wire             d1_nios_system_clock_4_in_end_xfer;
  wire             d1_nios_system_clock_5_in_end_xfer;
  wire             d1_nios_system_clock_6_in_end_xfer;
  wire             d1_nios_system_clock_7_in_end_xfer;
  wire             d1_nios_system_clock_8_in_end_xfer;
  wire             d1_nios_system_clock_9_in_end_xfer;
  wire             d1_onchip_memory2_0_s1_end_xfer;
  wire             d1_onchip_memory2_1_s1_end_xfer;
  wire             d1_onchip_memory2_2_s1_end_xfer;
  wire             d1_onchip_memory2_3_s1_end_xfer;
  wire             d1_performance_counter_0_control_slave_end_xfer;
  wire             d1_sdram_0_s1_end_xfer;
  wire             d1_sram_0_avalon_sram_slave_end_xfer;
  wire             d1_sysid_control_slave_end_xfer;
  wire             d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer;
  wire             jtag_uart_0_avalon_jtag_slave_address;
  wire             jtag_uart_0_avalon_jtag_slave_chipselect;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_irq;
  wire             jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_reset_n;
  wire             jtag_uart_0_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_writedata;
  wire             jtag_uart_1_avalon_jtag_slave_address;
  wire             jtag_uart_1_avalon_jtag_slave_chipselect;
  wire             jtag_uart_1_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_1_avalon_jtag_slave_irq;
  wire             jtag_uart_1_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_1_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_1_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_1_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_1_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_1_avalon_jtag_slave_reset_n;
  wire             jtag_uart_1_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_1_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_1_avalon_jtag_slave_writedata;
  wire             jtag_uart_2_avalon_jtag_slave_address;
  wire             jtag_uart_2_avalon_jtag_slave_chipselect;
  wire             jtag_uart_2_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_2_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_2_avalon_jtag_slave_irq;
  wire             jtag_uart_2_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_2_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_2_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_2_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_2_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_2_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_2_avalon_jtag_slave_reset_n;
  wire             jtag_uart_2_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_2_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_2_avalon_jtag_slave_writedata;
  wire             jtag_uart_3_avalon_jtag_slave_address;
  wire             jtag_uart_3_avalon_jtag_slave_chipselect;
  wire             jtag_uart_3_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_3_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_3_avalon_jtag_slave_irq;
  wire             jtag_uart_3_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_3_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_3_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_3_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_3_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_3_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_3_avalon_jtag_slave_reset_n;
  wire             jtag_uart_3_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_3_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_3_avalon_jtag_slave_writedata;
  wire    [  1: 0] keys_s1_address;
  wire             keys_s1_chipselect;
  wire    [ 31: 0] keys_s1_readdata;
  wire    [ 31: 0] keys_s1_readdata_from_sa;
  wire             keys_s1_reset_n;
  wire             keys_s1_write_n;
  wire    [ 31: 0] keys_s1_writedata;
  wire    [  1: 0] mailbox_0_s1_address;
  wire             mailbox_0_s1_chipselect;
  wire             mailbox_0_s1_read;
  wire    [ 31: 0] mailbox_0_s1_readdata;
  wire    [ 31: 0] mailbox_0_s1_readdata_from_sa;
  wire             mailbox_0_s1_reset_n;
  wire             mailbox_0_s1_write;
  wire    [ 31: 0] mailbox_0_s1_writedata;
  wire    [  1: 0] mailbox_1_s1_address;
  wire             mailbox_1_s1_chipselect;
  wire             mailbox_1_s1_read;
  wire    [ 31: 0] mailbox_1_s1_readdata;
  wire    [ 31: 0] mailbox_1_s1_readdata_from_sa;
  wire             mailbox_1_s1_reset_n;
  wire             mailbox_1_s1_write;
  wire    [ 31: 0] mailbox_1_s1_writedata;
  wire    [  1: 0] mailbox_2_s1_address;
  wire             mailbox_2_s1_chipselect;
  wire             mailbox_2_s1_read;
  wire    [ 31: 0] mailbox_2_s1_readdata;
  wire    [ 31: 0] mailbox_2_s1_readdata_from_sa;
  wire             mailbox_2_s1_reset_n;
  wire             mailbox_2_s1_write;
  wire    [ 31: 0] mailbox_2_s1_writedata;
  wire    [  1: 0] mailbox_3_s1_address;
  wire             mailbox_3_s1_chipselect;
  wire             mailbox_3_s1_read;
  wire    [ 31: 0] mailbox_3_s1_readdata;
  wire    [ 31: 0] mailbox_3_s1_readdata_from_sa;
  wire             mailbox_3_s1_reset_n;
  wire             mailbox_3_s1_write;
  wire    [ 31: 0] mailbox_3_s1_writedata;
  wire    [ 22: 0] nios_system_clock_0_in_address;
  wire    [  1: 0] nios_system_clock_0_in_byteenable;
  wire             nios_system_clock_0_in_endofpacket;
  wire             nios_system_clock_0_in_endofpacket_from_sa;
  wire    [ 21: 0] nios_system_clock_0_in_nativeaddress;
  wire             nios_system_clock_0_in_read;
  wire    [ 15: 0] nios_system_clock_0_in_readdata;
  wire    [ 15: 0] nios_system_clock_0_in_readdata_from_sa;
  wire             nios_system_clock_0_in_reset_n;
  wire             nios_system_clock_0_in_waitrequest;
  wire             nios_system_clock_0_in_waitrequest_from_sa;
  wire             nios_system_clock_0_in_write;
  wire    [ 15: 0] nios_system_clock_0_in_writedata;
  wire    [ 22: 0] nios_system_clock_0_out_address;
  wire    [ 22: 0] nios_system_clock_0_out_address_to_slave;
  wire    [  1: 0] nios_system_clock_0_out_byteenable;
  wire             nios_system_clock_0_out_endofpacket;
  wire             nios_system_clock_0_out_granted_sdram_0_s1;
  wire    [ 21: 0] nios_system_clock_0_out_nativeaddress;
  wire             nios_system_clock_0_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_0_out_read;
  wire             nios_system_clock_0_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register;
  wire    [ 15: 0] nios_system_clock_0_out_readdata;
  wire             nios_system_clock_0_out_requests_sdram_0_s1;
  wire             nios_system_clock_0_out_reset_n;
  wire             nios_system_clock_0_out_waitrequest;
  wire             nios_system_clock_0_out_write;
  wire    [ 15: 0] nios_system_clock_0_out_writedata;
  wire             nios_system_clock_10_in_address;
  wire             nios_system_clock_10_in_endofpacket;
  wire             nios_system_clock_10_in_endofpacket_from_sa;
  wire             nios_system_clock_10_in_nativeaddress;
  wire             nios_system_clock_10_in_read;
  wire    [  7: 0] nios_system_clock_10_in_readdata;
  wire    [  7: 0] nios_system_clock_10_in_readdata_from_sa;
  wire             nios_system_clock_10_in_reset_n;
  wire             nios_system_clock_10_in_waitrequest;
  wire             nios_system_clock_10_in_waitrequest_from_sa;
  wire             nios_system_clock_10_in_write;
  wire    [  7: 0] nios_system_clock_10_in_writedata;
  wire             nios_system_clock_10_out_address;
  wire             nios_system_clock_10_out_address_to_slave;
  wire             nios_system_clock_10_out_endofpacket;
  wire             nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_10_out_nativeaddress;
  wire             nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_10_out_read;
  wire             nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave;
  wire    [  7: 0] nios_system_clock_10_out_readdata;
  wire             nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_10_out_reset_n;
  wire             nios_system_clock_10_out_waitrequest;
  wire             nios_system_clock_10_out_write;
  wire    [  7: 0] nios_system_clock_10_out_writedata;
  wire             nios_system_clock_11_in_address;
  wire             nios_system_clock_11_in_endofpacket;
  wire             nios_system_clock_11_in_endofpacket_from_sa;
  wire             nios_system_clock_11_in_nativeaddress;
  wire             nios_system_clock_11_in_read;
  wire    [  7: 0] nios_system_clock_11_in_readdata;
  wire    [  7: 0] nios_system_clock_11_in_readdata_from_sa;
  wire             nios_system_clock_11_in_reset_n;
  wire             nios_system_clock_11_in_waitrequest;
  wire             nios_system_clock_11_in_waitrequest_from_sa;
  wire             nios_system_clock_11_in_write;
  wire    [  7: 0] nios_system_clock_11_in_writedata;
  wire             nios_system_clock_11_out_address;
  wire             nios_system_clock_11_out_address_to_slave;
  wire             nios_system_clock_11_out_endofpacket;
  wire             nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_11_out_nativeaddress;
  wire             nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_11_out_read;
  wire             nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave;
  wire    [  7: 0] nios_system_clock_11_out_readdata;
  wire             nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_11_out_reset_n;
  wire             nios_system_clock_11_out_waitrequest;
  wire             nios_system_clock_11_out_write;
  wire    [  7: 0] nios_system_clock_11_out_writedata;
  wire    [ 22: 0] nios_system_clock_1_in_address;
  wire    [  1: 0] nios_system_clock_1_in_byteenable;
  wire             nios_system_clock_1_in_endofpacket;
  wire             nios_system_clock_1_in_endofpacket_from_sa;
  wire    [ 21: 0] nios_system_clock_1_in_nativeaddress;
  wire             nios_system_clock_1_in_read;
  wire    [ 15: 0] nios_system_clock_1_in_readdata;
  wire    [ 15: 0] nios_system_clock_1_in_readdata_from_sa;
  wire             nios_system_clock_1_in_reset_n;
  wire             nios_system_clock_1_in_waitrequest;
  wire             nios_system_clock_1_in_waitrequest_from_sa;
  wire             nios_system_clock_1_in_write;
  wire    [ 15: 0] nios_system_clock_1_in_writedata;
  wire    [ 22: 0] nios_system_clock_1_out_address;
  wire    [ 22: 0] nios_system_clock_1_out_address_to_slave;
  wire    [  1: 0] nios_system_clock_1_out_byteenable;
  wire             nios_system_clock_1_out_endofpacket;
  wire             nios_system_clock_1_out_granted_sdram_0_s1;
  wire    [ 21: 0] nios_system_clock_1_out_nativeaddress;
  wire             nios_system_clock_1_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_1_out_read;
  wire             nios_system_clock_1_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register;
  wire    [ 15: 0] nios_system_clock_1_out_readdata;
  wire             nios_system_clock_1_out_requests_sdram_0_s1;
  wire             nios_system_clock_1_out_reset_n;
  wire             nios_system_clock_1_out_waitrequest;
  wire             nios_system_clock_1_out_write;
  wire    [ 15: 0] nios_system_clock_1_out_writedata;
  wire    [ 22: 0] nios_system_clock_2_in_address;
  wire    [  1: 0] nios_system_clock_2_in_byteenable;
  wire             nios_system_clock_2_in_endofpacket;
  wire             nios_system_clock_2_in_endofpacket_from_sa;
  wire    [ 21: 0] nios_system_clock_2_in_nativeaddress;
  wire             nios_system_clock_2_in_read;
  wire    [ 15: 0] nios_system_clock_2_in_readdata;
  wire    [ 15: 0] nios_system_clock_2_in_readdata_from_sa;
  wire             nios_system_clock_2_in_reset_n;
  wire             nios_system_clock_2_in_waitrequest;
  wire             nios_system_clock_2_in_waitrequest_from_sa;
  wire             nios_system_clock_2_in_write;
  wire    [ 15: 0] nios_system_clock_2_in_writedata;
  wire    [ 22: 0] nios_system_clock_2_out_address;
  wire    [ 22: 0] nios_system_clock_2_out_address_to_slave;
  wire    [  1: 0] nios_system_clock_2_out_byteenable;
  wire             nios_system_clock_2_out_endofpacket;
  wire             nios_system_clock_2_out_granted_sdram_0_s1;
  wire    [ 21: 0] nios_system_clock_2_out_nativeaddress;
  wire             nios_system_clock_2_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_2_out_read;
  wire             nios_system_clock_2_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register;
  wire    [ 15: 0] nios_system_clock_2_out_readdata;
  wire             nios_system_clock_2_out_requests_sdram_0_s1;
  wire             nios_system_clock_2_out_reset_n;
  wire             nios_system_clock_2_out_waitrequest;
  wire             nios_system_clock_2_out_write;
  wire    [ 15: 0] nios_system_clock_2_out_writedata;
  wire    [ 22: 0] nios_system_clock_3_in_address;
  wire    [  1: 0] nios_system_clock_3_in_byteenable;
  wire             nios_system_clock_3_in_endofpacket;
  wire             nios_system_clock_3_in_endofpacket_from_sa;
  wire    [ 21: 0] nios_system_clock_3_in_nativeaddress;
  wire             nios_system_clock_3_in_read;
  wire    [ 15: 0] nios_system_clock_3_in_readdata;
  wire    [ 15: 0] nios_system_clock_3_in_readdata_from_sa;
  wire             nios_system_clock_3_in_reset_n;
  wire             nios_system_clock_3_in_waitrequest;
  wire             nios_system_clock_3_in_waitrequest_from_sa;
  wire             nios_system_clock_3_in_write;
  wire    [ 15: 0] nios_system_clock_3_in_writedata;
  wire    [ 22: 0] nios_system_clock_3_out_address;
  wire    [ 22: 0] nios_system_clock_3_out_address_to_slave;
  wire    [  1: 0] nios_system_clock_3_out_byteenable;
  wire             nios_system_clock_3_out_endofpacket;
  wire             nios_system_clock_3_out_granted_sdram_0_s1;
  wire    [ 21: 0] nios_system_clock_3_out_nativeaddress;
  wire             nios_system_clock_3_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_3_out_read;
  wire             nios_system_clock_3_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register;
  wire    [ 15: 0] nios_system_clock_3_out_readdata;
  wire             nios_system_clock_3_out_requests_sdram_0_s1;
  wire             nios_system_clock_3_out_reset_n;
  wire             nios_system_clock_3_out_waitrequest;
  wire             nios_system_clock_3_out_write;
  wire    [ 15: 0] nios_system_clock_3_out_writedata;
  wire    [ 22: 0] nios_system_clock_4_in_address;
  wire    [  1: 0] nios_system_clock_4_in_byteenable;
  wire             nios_system_clock_4_in_endofpacket;
  wire             nios_system_clock_4_in_endofpacket_from_sa;
  wire    [ 21: 0] nios_system_clock_4_in_nativeaddress;
  wire             nios_system_clock_4_in_read;
  wire    [ 15: 0] nios_system_clock_4_in_readdata;
  wire    [ 15: 0] nios_system_clock_4_in_readdata_from_sa;
  wire             nios_system_clock_4_in_reset_n;
  wire             nios_system_clock_4_in_waitrequest;
  wire             nios_system_clock_4_in_waitrequest_from_sa;
  wire             nios_system_clock_4_in_write;
  wire    [ 15: 0] nios_system_clock_4_in_writedata;
  wire    [ 22: 0] nios_system_clock_4_out_address;
  wire    [ 22: 0] nios_system_clock_4_out_address_to_slave;
  wire    [  1: 0] nios_system_clock_4_out_byteenable;
  wire             nios_system_clock_4_out_endofpacket;
  wire             nios_system_clock_4_out_granted_sdram_0_s1;
  wire    [ 21: 0] nios_system_clock_4_out_nativeaddress;
  wire             nios_system_clock_4_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_4_out_read;
  wire             nios_system_clock_4_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register;
  wire    [ 15: 0] nios_system_clock_4_out_readdata;
  wire             nios_system_clock_4_out_requests_sdram_0_s1;
  wire             nios_system_clock_4_out_reset_n;
  wire             nios_system_clock_4_out_waitrequest;
  wire             nios_system_clock_4_out_write;
  wire    [ 15: 0] nios_system_clock_4_out_writedata;
  wire    [ 22: 0] nios_system_clock_5_in_address;
  wire    [  1: 0] nios_system_clock_5_in_byteenable;
  wire             nios_system_clock_5_in_endofpacket;
  wire             nios_system_clock_5_in_endofpacket_from_sa;
  wire    [ 21: 0] nios_system_clock_5_in_nativeaddress;
  wire             nios_system_clock_5_in_read;
  wire    [ 15: 0] nios_system_clock_5_in_readdata;
  wire    [ 15: 0] nios_system_clock_5_in_readdata_from_sa;
  wire             nios_system_clock_5_in_reset_n;
  wire             nios_system_clock_5_in_waitrequest;
  wire             nios_system_clock_5_in_waitrequest_from_sa;
  wire             nios_system_clock_5_in_write;
  wire    [ 15: 0] nios_system_clock_5_in_writedata;
  wire    [ 22: 0] nios_system_clock_5_out_address;
  wire    [ 22: 0] nios_system_clock_5_out_address_to_slave;
  wire    [  1: 0] nios_system_clock_5_out_byteenable;
  wire             nios_system_clock_5_out_endofpacket;
  wire             nios_system_clock_5_out_granted_sdram_0_s1;
  wire    [ 21: 0] nios_system_clock_5_out_nativeaddress;
  wire             nios_system_clock_5_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_5_out_read;
  wire             nios_system_clock_5_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register;
  wire    [ 15: 0] nios_system_clock_5_out_readdata;
  wire             nios_system_clock_5_out_requests_sdram_0_s1;
  wire             nios_system_clock_5_out_reset_n;
  wire             nios_system_clock_5_out_waitrequest;
  wire             nios_system_clock_5_out_write;
  wire    [ 15: 0] nios_system_clock_5_out_writedata;
  wire    [ 22: 0] nios_system_clock_6_in_address;
  wire    [  1: 0] nios_system_clock_6_in_byteenable;
  wire             nios_system_clock_6_in_endofpacket;
  wire             nios_system_clock_6_in_endofpacket_from_sa;
  wire    [ 21: 0] nios_system_clock_6_in_nativeaddress;
  wire             nios_system_clock_6_in_read;
  wire    [ 15: 0] nios_system_clock_6_in_readdata;
  wire    [ 15: 0] nios_system_clock_6_in_readdata_from_sa;
  wire             nios_system_clock_6_in_reset_n;
  wire             nios_system_clock_6_in_waitrequest;
  wire             nios_system_clock_6_in_waitrequest_from_sa;
  wire             nios_system_clock_6_in_write;
  wire    [ 15: 0] nios_system_clock_6_in_writedata;
  wire    [ 22: 0] nios_system_clock_6_out_address;
  wire    [ 22: 0] nios_system_clock_6_out_address_to_slave;
  wire    [  1: 0] nios_system_clock_6_out_byteenable;
  wire             nios_system_clock_6_out_endofpacket;
  wire             nios_system_clock_6_out_granted_sdram_0_s1;
  wire    [ 21: 0] nios_system_clock_6_out_nativeaddress;
  wire             nios_system_clock_6_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_6_out_read;
  wire             nios_system_clock_6_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register;
  wire    [ 15: 0] nios_system_clock_6_out_readdata;
  wire             nios_system_clock_6_out_requests_sdram_0_s1;
  wire             nios_system_clock_6_out_reset_n;
  wire             nios_system_clock_6_out_waitrequest;
  wire             nios_system_clock_6_out_write;
  wire    [ 15: 0] nios_system_clock_6_out_writedata;
  wire    [ 22: 0] nios_system_clock_7_in_address;
  wire    [  1: 0] nios_system_clock_7_in_byteenable;
  wire             nios_system_clock_7_in_endofpacket;
  wire             nios_system_clock_7_in_endofpacket_from_sa;
  wire    [ 21: 0] nios_system_clock_7_in_nativeaddress;
  wire             nios_system_clock_7_in_read;
  wire    [ 15: 0] nios_system_clock_7_in_readdata;
  wire    [ 15: 0] nios_system_clock_7_in_readdata_from_sa;
  wire             nios_system_clock_7_in_reset_n;
  wire             nios_system_clock_7_in_waitrequest;
  wire             nios_system_clock_7_in_waitrequest_from_sa;
  wire             nios_system_clock_7_in_write;
  wire    [ 15: 0] nios_system_clock_7_in_writedata;
  wire    [ 22: 0] nios_system_clock_7_out_address;
  wire    [ 22: 0] nios_system_clock_7_out_address_to_slave;
  wire    [  1: 0] nios_system_clock_7_out_byteenable;
  wire             nios_system_clock_7_out_endofpacket;
  wire             nios_system_clock_7_out_granted_sdram_0_s1;
  wire    [ 21: 0] nios_system_clock_7_out_nativeaddress;
  wire             nios_system_clock_7_out_qualified_request_sdram_0_s1;
  wire             nios_system_clock_7_out_read;
  wire             nios_system_clock_7_out_read_data_valid_sdram_0_s1;
  wire             nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register;
  wire    [ 15: 0] nios_system_clock_7_out_readdata;
  wire             nios_system_clock_7_out_requests_sdram_0_s1;
  wire             nios_system_clock_7_out_reset_n;
  wire             nios_system_clock_7_out_waitrequest;
  wire             nios_system_clock_7_out_write;
  wire    [ 15: 0] nios_system_clock_7_out_writedata;
  wire             nios_system_clock_8_in_address;
  wire             nios_system_clock_8_in_endofpacket;
  wire             nios_system_clock_8_in_endofpacket_from_sa;
  wire             nios_system_clock_8_in_nativeaddress;
  wire             nios_system_clock_8_in_read;
  wire    [  7: 0] nios_system_clock_8_in_readdata;
  wire    [  7: 0] nios_system_clock_8_in_readdata_from_sa;
  wire             nios_system_clock_8_in_reset_n;
  wire             nios_system_clock_8_in_waitrequest;
  wire             nios_system_clock_8_in_waitrequest_from_sa;
  wire             nios_system_clock_8_in_write;
  wire    [  7: 0] nios_system_clock_8_in_writedata;
  wire             nios_system_clock_8_out_address;
  wire             nios_system_clock_8_out_address_to_slave;
  wire             nios_system_clock_8_out_endofpacket;
  wire             nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_8_out_nativeaddress;
  wire             nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_8_out_read;
  wire             nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave;
  wire    [  7: 0] nios_system_clock_8_out_readdata;
  wire             nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_8_out_reset_n;
  wire             nios_system_clock_8_out_waitrequest;
  wire             nios_system_clock_8_out_write;
  wire    [  7: 0] nios_system_clock_8_out_writedata;
  wire             nios_system_clock_9_in_address;
  wire             nios_system_clock_9_in_endofpacket;
  wire             nios_system_clock_9_in_endofpacket_from_sa;
  wire             nios_system_clock_9_in_nativeaddress;
  wire             nios_system_clock_9_in_read;
  wire    [  7: 0] nios_system_clock_9_in_readdata;
  wire    [  7: 0] nios_system_clock_9_in_readdata_from_sa;
  wire             nios_system_clock_9_in_reset_n;
  wire             nios_system_clock_9_in_waitrequest;
  wire             nios_system_clock_9_in_waitrequest_from_sa;
  wire             nios_system_clock_9_in_write;
  wire    [  7: 0] nios_system_clock_9_in_writedata;
  wire             nios_system_clock_9_out_address;
  wire             nios_system_clock_9_out_address_to_slave;
  wire             nios_system_clock_9_out_endofpacket;
  wire             nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_9_out_nativeaddress;
  wire             nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_9_out_read;
  wire             nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave;
  wire    [  7: 0] nios_system_clock_9_out_readdata;
  wire             nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave;
  wire             nios_system_clock_9_out_reset_n;
  wire             nios_system_clock_9_out_waitrequest;
  wire             nios_system_clock_9_out_write;
  wire    [  7: 0] nios_system_clock_9_out_writedata;
  wire    [  6: 0] onchip_memory2_0_s1_address;
  wire    [  3: 0] onchip_memory2_0_s1_byteenable;
  wire             onchip_memory2_0_s1_chipselect;
  wire             onchip_memory2_0_s1_clken;
  wire    [ 31: 0] onchip_memory2_0_s1_readdata;
  wire    [ 31: 0] onchip_memory2_0_s1_readdata_from_sa;
  wire             onchip_memory2_0_s1_reset;
  wire             onchip_memory2_0_s1_write;
  wire    [ 31: 0] onchip_memory2_0_s1_writedata;
  wire    [  6: 0] onchip_memory2_1_s1_address;
  wire    [  3: 0] onchip_memory2_1_s1_byteenable;
  wire             onchip_memory2_1_s1_chipselect;
  wire             onchip_memory2_1_s1_clken;
  wire    [ 31: 0] onchip_memory2_1_s1_readdata;
  wire    [ 31: 0] onchip_memory2_1_s1_readdata_from_sa;
  wire             onchip_memory2_1_s1_reset;
  wire             onchip_memory2_1_s1_write;
  wire    [ 31: 0] onchip_memory2_1_s1_writedata;
  wire    [  6: 0] onchip_memory2_2_s1_address;
  wire    [  3: 0] onchip_memory2_2_s1_byteenable;
  wire             onchip_memory2_2_s1_chipselect;
  wire             onchip_memory2_2_s1_clken;
  wire    [ 31: 0] onchip_memory2_2_s1_readdata;
  wire    [ 31: 0] onchip_memory2_2_s1_readdata_from_sa;
  wire             onchip_memory2_2_s1_reset;
  wire             onchip_memory2_2_s1_write;
  wire    [ 31: 0] onchip_memory2_2_s1_writedata;
  wire    [  6: 0] onchip_memory2_3_s1_address;
  wire    [  3: 0] onchip_memory2_3_s1_byteenable;
  wire             onchip_memory2_3_s1_chipselect;
  wire             onchip_memory2_3_s1_clken;
  wire    [ 31: 0] onchip_memory2_3_s1_readdata;
  wire    [ 31: 0] onchip_memory2_3_s1_readdata_from_sa;
  wire             onchip_memory2_3_s1_reset;
  wire             onchip_memory2_3_s1_write;
  wire    [ 31: 0] onchip_memory2_3_s1_writedata;
  wire             out_clk_clocks_0_SDRAM_CLK;
  wire             out_clk_clocks_0_VGA_CLK;
  wire             out_clk_clocks_0_sys_clk;
  wire    [  3: 0] performance_counter_0_control_slave_address;
  wire             performance_counter_0_control_slave_begintransfer;
  wire    [ 31: 0] performance_counter_0_control_slave_readdata;
  wire    [ 31: 0] performance_counter_0_control_slave_readdata_from_sa;
  wire             performance_counter_0_control_slave_reset_n;
  wire             performance_counter_0_control_slave_write;
  wire    [ 31: 0] performance_counter_0_control_slave_writedata;
  wire             reset_n_sources;
  wire    [ 21: 0] sdram_0_s1_address;
  wire    [  1: 0] sdram_0_s1_byteenable_n;
  wire             sdram_0_s1_chipselect;
  wire             sdram_0_s1_read_n;
  wire    [ 15: 0] sdram_0_s1_readdata;
  wire    [ 15: 0] sdram_0_s1_readdata_from_sa;
  wire             sdram_0_s1_readdatavalid;
  wire             sdram_0_s1_reset_n;
  wire             sdram_0_s1_waitrequest;
  wire             sdram_0_s1_waitrequest_from_sa;
  wire             sdram_0_s1_write_n;
  wire    [ 15: 0] sdram_0_s1_writedata;
  wire             sdram_clk;
  wire             sdram_clk_reset_n;
  wire    [ 17: 0] sram_0_avalon_sram_slave_address;
  wire    [  1: 0] sram_0_avalon_sram_slave_byteenable;
  wire             sram_0_avalon_sram_slave_read;
  wire    [ 15: 0] sram_0_avalon_sram_slave_readdata;
  wire    [ 15: 0] sram_0_avalon_sram_slave_readdata_from_sa;
  wire             sram_0_avalon_sram_slave_readdatavalid;
  wire             sram_0_avalon_sram_slave_reset;
  wire             sram_0_avalon_sram_slave_write;
  wire    [ 15: 0] sram_0_avalon_sram_slave_writedata;
  wire             sys_clk;
  wire             sys_clk_reset_n;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_clock;
  wire    [ 31: 0] sysid_control_slave_readdata;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  wire             sysid_control_slave_reset_n;
  wire             vga_clock;
  wire             vga_clock_reset_n;
  wire    [ 29: 0] video_dual_clock_buffer_0_avalon_dc_buffer_sink_data;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_sink_endofpacket;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_sink_startofpacket;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_sink_valid;
  wire    [ 29: 0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;
  wire             video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;
  wire    [  1: 0] video_pixel_buffer_dma_0_avalon_control_slave_address;
  wire    [  3: 0] video_pixel_buffer_dma_0_avalon_control_slave_byteenable;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_read;
  wire    [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_readdata;
  wire    [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa;
  wire             video_pixel_buffer_dma_0_avalon_control_slave_write;
  wire    [ 31: 0] video_pixel_buffer_dma_0_avalon_control_slave_writedata;
  wire    [ 31: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address;
  wire    [ 31: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock;
  wire    [  1: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_read;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave_shift_register;
  wire    [ 31: 0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_reset;
  wire             video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest;
  wire    [ 23: 0] video_pixel_buffer_dma_0_avalon_pixel_source_data;
  wire             video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket;
  wire             video_pixel_buffer_dma_0_avalon_pixel_source_ready;
  wire             video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket;
  wire             video_pixel_buffer_dma_0_avalon_pixel_source_valid;
  wire    [ 23: 0] video_rgb_resampler_0_avalon_rgb_sink_data;
  wire             video_rgb_resampler_0_avalon_rgb_sink_endofpacket;
  wire             video_rgb_resampler_0_avalon_rgb_sink_ready;
  wire             video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa;
  wire             video_rgb_resampler_0_avalon_rgb_sink_reset;
  wire             video_rgb_resampler_0_avalon_rgb_sink_startofpacket;
  wire             video_rgb_resampler_0_avalon_rgb_sink_valid;
  wire    [ 29: 0] video_rgb_resampler_0_avalon_rgb_source_data;
  wire             video_rgb_resampler_0_avalon_rgb_source_endofpacket;
  wire             video_rgb_resampler_0_avalon_rgb_source_ready;
  wire             video_rgb_resampler_0_avalon_rgb_source_startofpacket;
  wire             video_rgb_resampler_0_avalon_rgb_source_valid;
  wire    [ 29: 0] video_scaler_0_avalon_scaler_sink_data;
  wire             video_scaler_0_avalon_scaler_sink_endofpacket;
  wire             video_scaler_0_avalon_scaler_sink_ready;
  wire             video_scaler_0_avalon_scaler_sink_ready_from_sa;
  wire             video_scaler_0_avalon_scaler_sink_reset;
  wire             video_scaler_0_avalon_scaler_sink_startofpacket;
  wire             video_scaler_0_avalon_scaler_sink_valid;
  wire    [ 29: 0] video_scaler_0_avalon_scaler_source_data;
  wire             video_scaler_0_avalon_scaler_source_endofpacket;
  wire             video_scaler_0_avalon_scaler_source_ready;
  wire             video_scaler_0_avalon_scaler_source_startofpacket;
  wire             video_scaler_0_avalon_scaler_source_valid;
  wire    [ 29: 0] video_vga_controller_0_avalon_vga_sink_data;
  wire             video_vga_controller_0_avalon_vga_sink_endofpacket;
  wire             video_vga_controller_0_avalon_vga_sink_ready;
  wire             video_vga_controller_0_avalon_vga_sink_ready_from_sa;
  wire             video_vga_controller_0_avalon_vga_sink_reset;
  wire             video_vga_controller_0_avalon_vga_sink_startofpacket;
  wire             video_vga_controller_0_avalon_vga_sink_valid;
  wire    [ 11: 0] zs_addr_from_the_sdram_0;
  wire    [  1: 0] zs_ba_from_the_sdram_0;
  wire             zs_cas_n_from_the_sdram_0;
  wire             zs_cke_from_the_sdram_0;
  wire             zs_cs_n_from_the_sdram_0;
  wire    [ 15: 0] zs_dq_to_and_from_the_sdram_0;
  wire    [  1: 0] zs_dqm_from_the_sdram_0;
  wire             zs_ras_n_from_the_sdram_0;
  wire             zs_we_n_from_the_sdram_0;
  clocks_0_avalon_clocks_slave_arbitrator the_clocks_0_avalon_clocks_slave
    (
      .clk                                                                     (clk_0),
      .clocks_0_avalon_clocks_slave_address                                    (clocks_0_avalon_clocks_slave_address),
      .clocks_0_avalon_clocks_slave_readdata                                   (clocks_0_avalon_clocks_slave_readdata),
      .clocks_0_avalon_clocks_slave_readdata_from_sa                           (clocks_0_avalon_clocks_slave_readdata_from_sa),
      .d1_clocks_0_avalon_clocks_slave_end_xfer                                (d1_clocks_0_avalon_clocks_slave_end_xfer),
      .nios_system_clock_10_out_address_to_slave                               (nios_system_clock_10_out_address_to_slave),
      .nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave           (nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave),
      .nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave (nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave),
      .nios_system_clock_10_out_read                                           (nios_system_clock_10_out_read),
      .nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave   (nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave),
      .nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave          (nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave),
      .nios_system_clock_10_out_write                                          (nios_system_clock_10_out_write),
      .nios_system_clock_11_out_address_to_slave                               (nios_system_clock_11_out_address_to_slave),
      .nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave           (nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave),
      .nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave (nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave),
      .nios_system_clock_11_out_read                                           (nios_system_clock_11_out_read),
      .nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave   (nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave),
      .nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave          (nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave),
      .nios_system_clock_11_out_write                                          (nios_system_clock_11_out_write),
      .nios_system_clock_8_out_address_to_slave                                (nios_system_clock_8_out_address_to_slave),
      .nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave            (nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave),
      .nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave  (nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave),
      .nios_system_clock_8_out_read                                            (nios_system_clock_8_out_read),
      .nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave    (nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave),
      .nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave           (nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave),
      .nios_system_clock_8_out_write                                           (nios_system_clock_8_out_write),
      .nios_system_clock_9_out_address_to_slave                                (nios_system_clock_9_out_address_to_slave),
      .nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave            (nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave),
      .nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave  (nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave),
      .nios_system_clock_9_out_read                                            (nios_system_clock_9_out_read),
      .nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave    (nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave),
      .nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave           (nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave),
      .nios_system_clock_9_out_write                                           (nios_system_clock_9_out_write),
      .reset_n                                                                 (clk_0_reset_n)
    );

  //sdram_clk out_clk assignment, which is an e_assign
  assign sdram_clk = out_clk_clocks_0_SDRAM_CLK;

  //vga_clock out_clk assignment, which is an e_assign
  assign vga_clock = out_clk_clocks_0_VGA_CLK;

  //sys_clk out_clk assignment, which is an e_assign
  assign sys_clk = out_clk_clocks_0_sys_clk;

  clocks_0 the_clocks_0
    (
      .CLOCK_50  (clk_0),
      .SDRAM_CLK (out_clk_clocks_0_SDRAM_CLK),
      .VGA_CLK   (out_clk_clocks_0_VGA_CLK),
      .address   (clocks_0_avalon_clocks_slave_address),
      .readdata  (clocks_0_avalon_clocks_slave_readdata),
      .sys_clk   (out_clk_clocks_0_sys_clk)
    );

  cpu_0_jtag_debug_module_arbitrator the_cpu_0_jtag_debug_module
    (
      .clk                                                                       (sys_clk),
      .cpu_0_data_master_address_to_slave                                        (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                              (cpu_0_data_master_byteenable),
      .cpu_0_data_master_debugaccess                                             (cpu_0_data_master_debugaccess),
      .cpu_0_data_master_granted_cpu_0_jtag_debug_module                         (cpu_0_data_master_granted_cpu_0_jtag_debug_module),
      .cpu_0_data_master_latency_counter                                         (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module               (cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module),
      .cpu_0_data_master_read                                                    (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module                 (cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_cpu_0_jtag_debug_module                        (cpu_0_data_master_requests_cpu_0_jtag_debug_module),
      .cpu_0_data_master_write                                                   (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                               (cpu_0_data_master_writedata),
      .cpu_0_instruction_master_address_to_slave                                 (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_granted_cpu_0_jtag_debug_module                  (cpu_0_instruction_master_granted_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_latency_counter                                  (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module        (cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_read                                             (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module          (cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_requests_cpu_0_jtag_debug_module                 (cpu_0_instruction_master_requests_cpu_0_jtag_debug_module),
      .cpu_0_jtag_debug_module_address                                           (cpu_0_jtag_debug_module_address),
      .cpu_0_jtag_debug_module_begintransfer                                     (cpu_0_jtag_debug_module_begintransfer),
      .cpu_0_jtag_debug_module_byteenable                                        (cpu_0_jtag_debug_module_byteenable),
      .cpu_0_jtag_debug_module_chipselect                                        (cpu_0_jtag_debug_module_chipselect),
      .cpu_0_jtag_debug_module_debugaccess                                       (cpu_0_jtag_debug_module_debugaccess),
      .cpu_0_jtag_debug_module_readdata                                          (cpu_0_jtag_debug_module_readdata),
      .cpu_0_jtag_debug_module_readdata_from_sa                                  (cpu_0_jtag_debug_module_readdata_from_sa),
      .cpu_0_jtag_debug_module_resetrequest                                      (cpu_0_jtag_debug_module_resetrequest),
      .cpu_0_jtag_debug_module_resetrequest_from_sa                              (cpu_0_jtag_debug_module_resetrequest_from_sa),
      .cpu_0_jtag_debug_module_write                                             (cpu_0_jtag_debug_module_write),
      .cpu_0_jtag_debug_module_writedata                                         (cpu_0_jtag_debug_module_writedata),
      .d1_cpu_0_jtag_debug_module_end_xfer                                       (d1_cpu_0_jtag_debug_module_end_xfer),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  cpu_0_custom_instruction_master_arbitrator the_cpu_0_custom_instruction_master
    (
      .clk                                                                                         (sys_clk),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa                          (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa                        (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select                                (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select),
      .cpu_0_custom_instruction_master_multi_done                                                  (cpu_0_custom_instruction_master_multi_done),
      .cpu_0_custom_instruction_master_multi_result                                                (cpu_0_custom_instruction_master_multi_result),
      .cpu_0_custom_instruction_master_multi_start                                                 (cpu_0_custom_instruction_master_multi_start),
      .cpu_0_custom_instruction_master_reset_n                                                     (cpu_0_custom_instruction_master_reset_n),
      .cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1 (cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1),
      .reset_n                                                                                     (sys_clk_reset_n)
    );

  cpu_0_data_master_arbitrator the_cpu_0_data_master
    (
      .clk                                                                               (sys_clk),
      .cpu_0_data_master_address                                                         (cpu_0_data_master_address),
      .cpu_0_data_master_address_to_slave                                                (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                                      (cpu_0_data_master_byteenable),
      .cpu_0_data_master_byteenable_nios_system_clock_3_in                               (cpu_0_data_master_byteenable_nios_system_clock_3_in),
      .cpu_0_data_master_byteenable_nios_system_clock_9_in                               (cpu_0_data_master_byteenable_nios_system_clock_9_in),
      .cpu_0_data_master_byteenable_sram_0_avalon_sram_slave                             (cpu_0_data_master_byteenable_sram_0_avalon_sram_slave),
      .cpu_0_data_master_dbs_address                                                     (cpu_0_data_master_dbs_address),
      .cpu_0_data_master_dbs_write_16                                                    (cpu_0_data_master_dbs_write_16),
      .cpu_0_data_master_dbs_write_8                                                     (cpu_0_data_master_dbs_write_8),
      .cpu_0_data_master_granted_cpu_0_jtag_debug_module                                 (cpu_0_data_master_granted_cpu_0_jtag_debug_module),
      .cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave                           (cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_granted_keys_s1                                                 (cpu_0_data_master_granted_keys_s1),
      .cpu_0_data_master_granted_mailbox_0_s1                                            (cpu_0_data_master_granted_mailbox_0_s1),
      .cpu_0_data_master_granted_mailbox_1_s1                                            (cpu_0_data_master_granted_mailbox_1_s1),
      .cpu_0_data_master_granted_mailbox_2_s1                                            (cpu_0_data_master_granted_mailbox_2_s1),
      .cpu_0_data_master_granted_mailbox_3_s1                                            (cpu_0_data_master_granted_mailbox_3_s1),
      .cpu_0_data_master_granted_nios_system_clock_3_in                                  (cpu_0_data_master_granted_nios_system_clock_3_in),
      .cpu_0_data_master_granted_nios_system_clock_9_in                                  (cpu_0_data_master_granted_nios_system_clock_9_in),
      .cpu_0_data_master_granted_onchip_memory2_0_s1                                     (cpu_0_data_master_granted_onchip_memory2_0_s1),
      .cpu_0_data_master_granted_onchip_memory2_1_s1                                     (cpu_0_data_master_granted_onchip_memory2_1_s1),
      .cpu_0_data_master_granted_onchip_memory2_2_s1                                     (cpu_0_data_master_granted_onchip_memory2_2_s1),
      .cpu_0_data_master_granted_onchip_memory2_3_s1                                     (cpu_0_data_master_granted_onchip_memory2_3_s1),
      .cpu_0_data_master_granted_performance_counter_0_control_slave                     (cpu_0_data_master_granted_performance_counter_0_control_slave),
      .cpu_0_data_master_granted_sram_0_avalon_sram_slave                                (cpu_0_data_master_granted_sram_0_avalon_sram_slave),
      .cpu_0_data_master_granted_sysid_control_slave                                     (cpu_0_data_master_granted_sysid_control_slave),
      .cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave           (cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_0_data_master_irq                                                             (cpu_0_data_master_irq),
      .cpu_0_data_master_latency_counter                                                 (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module                       (cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module),
      .cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave                 (cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_qualified_request_keys_s1                                       (cpu_0_data_master_qualified_request_keys_s1),
      .cpu_0_data_master_qualified_request_mailbox_0_s1                                  (cpu_0_data_master_qualified_request_mailbox_0_s1),
      .cpu_0_data_master_qualified_request_mailbox_1_s1                                  (cpu_0_data_master_qualified_request_mailbox_1_s1),
      .cpu_0_data_master_qualified_request_mailbox_2_s1                                  (cpu_0_data_master_qualified_request_mailbox_2_s1),
      .cpu_0_data_master_qualified_request_mailbox_3_s1                                  (cpu_0_data_master_qualified_request_mailbox_3_s1),
      .cpu_0_data_master_qualified_request_nios_system_clock_3_in                        (cpu_0_data_master_qualified_request_nios_system_clock_3_in),
      .cpu_0_data_master_qualified_request_nios_system_clock_9_in                        (cpu_0_data_master_qualified_request_nios_system_clock_9_in),
      .cpu_0_data_master_qualified_request_onchip_memory2_0_s1                           (cpu_0_data_master_qualified_request_onchip_memory2_0_s1),
      .cpu_0_data_master_qualified_request_onchip_memory2_1_s1                           (cpu_0_data_master_qualified_request_onchip_memory2_1_s1),
      .cpu_0_data_master_qualified_request_onchip_memory2_2_s1                           (cpu_0_data_master_qualified_request_onchip_memory2_2_s1),
      .cpu_0_data_master_qualified_request_onchip_memory2_3_s1                           (cpu_0_data_master_qualified_request_onchip_memory2_3_s1),
      .cpu_0_data_master_qualified_request_performance_counter_0_control_slave           (cpu_0_data_master_qualified_request_performance_counter_0_control_slave),
      .cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave                      (cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_0_data_master_qualified_request_sysid_control_slave                           (cpu_0_data_master_qualified_request_sysid_control_slave),
      .cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave (cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_0_data_master_read                                                            (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module                         (cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module),
      .cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave                   (cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_read_data_valid_keys_s1                                         (cpu_0_data_master_read_data_valid_keys_s1),
      .cpu_0_data_master_read_data_valid_mailbox_0_s1                                    (cpu_0_data_master_read_data_valid_mailbox_0_s1),
      .cpu_0_data_master_read_data_valid_mailbox_1_s1                                    (cpu_0_data_master_read_data_valid_mailbox_1_s1),
      .cpu_0_data_master_read_data_valid_mailbox_2_s1                                    (cpu_0_data_master_read_data_valid_mailbox_2_s1),
      .cpu_0_data_master_read_data_valid_mailbox_3_s1                                    (cpu_0_data_master_read_data_valid_mailbox_3_s1),
      .cpu_0_data_master_read_data_valid_nios_system_clock_3_in                          (cpu_0_data_master_read_data_valid_nios_system_clock_3_in),
      .cpu_0_data_master_read_data_valid_nios_system_clock_9_in                          (cpu_0_data_master_read_data_valid_nios_system_clock_9_in),
      .cpu_0_data_master_read_data_valid_onchip_memory2_0_s1                             (cpu_0_data_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_0_data_master_read_data_valid_onchip_memory2_1_s1                             (cpu_0_data_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_0_data_master_read_data_valid_onchip_memory2_2_s1                             (cpu_0_data_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_0_data_master_read_data_valid_onchip_memory2_3_s1                             (cpu_0_data_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_0_data_master_read_data_valid_performance_counter_0_control_slave             (cpu_0_data_master_read_data_valid_performance_counter_0_control_slave),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave                        (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register         (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_read_data_valid_sysid_control_slave                             (cpu_0_data_master_read_data_valid_sysid_control_slave),
      .cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave   (cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_0_data_master_readdata                                                        (cpu_0_data_master_readdata),
      .cpu_0_data_master_readdatavalid                                                   (cpu_0_data_master_readdatavalid),
      .cpu_0_data_master_requests_cpu_0_jtag_debug_module                                (cpu_0_data_master_requests_cpu_0_jtag_debug_module),
      .cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave                          (cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_requests_keys_s1                                                (cpu_0_data_master_requests_keys_s1),
      .cpu_0_data_master_requests_mailbox_0_s1                                           (cpu_0_data_master_requests_mailbox_0_s1),
      .cpu_0_data_master_requests_mailbox_1_s1                                           (cpu_0_data_master_requests_mailbox_1_s1),
      .cpu_0_data_master_requests_mailbox_2_s1                                           (cpu_0_data_master_requests_mailbox_2_s1),
      .cpu_0_data_master_requests_mailbox_3_s1                                           (cpu_0_data_master_requests_mailbox_3_s1),
      .cpu_0_data_master_requests_nios_system_clock_3_in                                 (cpu_0_data_master_requests_nios_system_clock_3_in),
      .cpu_0_data_master_requests_nios_system_clock_9_in                                 (cpu_0_data_master_requests_nios_system_clock_9_in),
      .cpu_0_data_master_requests_onchip_memory2_0_s1                                    (cpu_0_data_master_requests_onchip_memory2_0_s1),
      .cpu_0_data_master_requests_onchip_memory2_1_s1                                    (cpu_0_data_master_requests_onchip_memory2_1_s1),
      .cpu_0_data_master_requests_onchip_memory2_2_s1                                    (cpu_0_data_master_requests_onchip_memory2_2_s1),
      .cpu_0_data_master_requests_onchip_memory2_3_s1                                    (cpu_0_data_master_requests_onchip_memory2_3_s1),
      .cpu_0_data_master_requests_performance_counter_0_control_slave                    (cpu_0_data_master_requests_performance_counter_0_control_slave),
      .cpu_0_data_master_requests_sram_0_avalon_sram_slave                               (cpu_0_data_master_requests_sram_0_avalon_sram_slave),
      .cpu_0_data_master_requests_sysid_control_slave                                    (cpu_0_data_master_requests_sysid_control_slave),
      .cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave          (cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_0_data_master_waitrequest                                                     (cpu_0_data_master_waitrequest),
      .cpu_0_data_master_write                                                           (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                                       (cpu_0_data_master_writedata),
      .cpu_0_jtag_debug_module_readdata_from_sa                                          (cpu_0_jtag_debug_module_readdata_from_sa),
      .d1_cpu_0_jtag_debug_module_end_xfer                                               (d1_cpu_0_jtag_debug_module_end_xfer),
      .d1_jtag_uart_0_avalon_jtag_slave_end_xfer                                         (d1_jtag_uart_0_avalon_jtag_slave_end_xfer),
      .d1_keys_s1_end_xfer                                                               (d1_keys_s1_end_xfer),
      .d1_mailbox_0_s1_end_xfer                                                          (d1_mailbox_0_s1_end_xfer),
      .d1_mailbox_1_s1_end_xfer                                                          (d1_mailbox_1_s1_end_xfer),
      .d1_mailbox_2_s1_end_xfer                                                          (d1_mailbox_2_s1_end_xfer),
      .d1_mailbox_3_s1_end_xfer                                                          (d1_mailbox_3_s1_end_xfer),
      .d1_nios_system_clock_3_in_end_xfer                                                (d1_nios_system_clock_3_in_end_xfer),
      .d1_nios_system_clock_9_in_end_xfer                                                (d1_nios_system_clock_9_in_end_xfer),
      .d1_onchip_memory2_0_s1_end_xfer                                                   (d1_onchip_memory2_0_s1_end_xfer),
      .d1_onchip_memory2_1_s1_end_xfer                                                   (d1_onchip_memory2_1_s1_end_xfer),
      .d1_onchip_memory2_2_s1_end_xfer                                                   (d1_onchip_memory2_2_s1_end_xfer),
      .d1_onchip_memory2_3_s1_end_xfer                                                   (d1_onchip_memory2_3_s1_end_xfer),
      .d1_performance_counter_0_control_slave_end_xfer                                   (d1_performance_counter_0_control_slave_end_xfer),
      .d1_sram_0_avalon_sram_slave_end_xfer                                              (d1_sram_0_avalon_sram_slave_end_xfer),
      .d1_sysid_control_slave_end_xfer                                                   (d1_sysid_control_slave_end_xfer),
      .d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer                         (d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer),
      .jtag_uart_0_avalon_jtag_slave_irq_from_sa                                         (jtag_uart_0_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_0_avalon_jtag_slave_readdata_from_sa                                    (jtag_uart_0_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa                                 (jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa),
      .keys_s1_readdata_from_sa                                                          (keys_s1_readdata_from_sa),
      .mailbox_0_s1_readdata_from_sa                                                     (mailbox_0_s1_readdata_from_sa),
      .mailbox_1_s1_readdata_from_sa                                                     (mailbox_1_s1_readdata_from_sa),
      .mailbox_2_s1_readdata_from_sa                                                     (mailbox_2_s1_readdata_from_sa),
      .mailbox_3_s1_readdata_from_sa                                                     (mailbox_3_s1_readdata_from_sa),
      .nios_system_clock_3_in_readdata_from_sa                                           (nios_system_clock_3_in_readdata_from_sa),
      .nios_system_clock_3_in_waitrequest_from_sa                                        (nios_system_clock_3_in_waitrequest_from_sa),
      .nios_system_clock_9_in_readdata_from_sa                                           (nios_system_clock_9_in_readdata_from_sa),
      .nios_system_clock_9_in_waitrequest_from_sa                                        (nios_system_clock_9_in_waitrequest_from_sa),
      .onchip_memory2_0_s1_readdata_from_sa                                              (onchip_memory2_0_s1_readdata_from_sa),
      .onchip_memory2_1_s1_readdata_from_sa                                              (onchip_memory2_1_s1_readdata_from_sa),
      .onchip_memory2_2_s1_readdata_from_sa                                              (onchip_memory2_2_s1_readdata_from_sa),
      .onchip_memory2_3_s1_readdata_from_sa                                              (onchip_memory2_3_s1_readdata_from_sa),
      .performance_counter_0_control_slave_readdata_from_sa                              (performance_counter_0_control_slave_readdata_from_sa),
      .reset_n                                                                           (sys_clk_reset_n),
      .sram_0_avalon_sram_slave_readdata_from_sa                                         (sram_0_avalon_sram_slave_readdata_from_sa),
      .sysid_control_slave_readdata_from_sa                                              (sysid_control_slave_readdata_from_sa),
      .video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa                    (video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa)
    );

  cpu_0_instruction_master_arbitrator the_cpu_0_instruction_master
    (
      .clk                                                                (sys_clk),
      .cpu_0_instruction_master_address                                   (cpu_0_instruction_master_address),
      .cpu_0_instruction_master_address_to_slave                          (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_dbs_address                               (cpu_0_instruction_master_dbs_address),
      .cpu_0_instruction_master_granted_cpu_0_jtag_debug_module           (cpu_0_instruction_master_granted_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_granted_nios_system_clock_2_in            (cpu_0_instruction_master_granted_nios_system_clock_2_in),
      .cpu_0_instruction_master_granted_onchip_memory2_0_s1               (cpu_0_instruction_master_granted_onchip_memory2_0_s1),
      .cpu_0_instruction_master_granted_onchip_memory2_1_s1               (cpu_0_instruction_master_granted_onchip_memory2_1_s1),
      .cpu_0_instruction_master_granted_onchip_memory2_2_s1               (cpu_0_instruction_master_granted_onchip_memory2_2_s1),
      .cpu_0_instruction_master_granted_onchip_memory2_3_s1               (cpu_0_instruction_master_granted_onchip_memory2_3_s1),
      .cpu_0_instruction_master_latency_counter                           (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module (cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_qualified_request_nios_system_clock_2_in  (cpu_0_instruction_master_qualified_request_nios_system_clock_2_in),
      .cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1     (cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1),
      .cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1     (cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1),
      .cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1     (cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1),
      .cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1     (cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1),
      .cpu_0_instruction_master_read                                      (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module   (cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in    (cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in),
      .cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1       (cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1       (cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1       (cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1       (cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_0_instruction_master_readdata                                  (cpu_0_instruction_master_readdata),
      .cpu_0_instruction_master_readdatavalid                             (cpu_0_instruction_master_readdatavalid),
      .cpu_0_instruction_master_requests_cpu_0_jtag_debug_module          (cpu_0_instruction_master_requests_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_requests_nios_system_clock_2_in           (cpu_0_instruction_master_requests_nios_system_clock_2_in),
      .cpu_0_instruction_master_requests_onchip_memory2_0_s1              (cpu_0_instruction_master_requests_onchip_memory2_0_s1),
      .cpu_0_instruction_master_requests_onchip_memory2_1_s1              (cpu_0_instruction_master_requests_onchip_memory2_1_s1),
      .cpu_0_instruction_master_requests_onchip_memory2_2_s1              (cpu_0_instruction_master_requests_onchip_memory2_2_s1),
      .cpu_0_instruction_master_requests_onchip_memory2_3_s1              (cpu_0_instruction_master_requests_onchip_memory2_3_s1),
      .cpu_0_instruction_master_waitrequest                               (cpu_0_instruction_master_waitrequest),
      .cpu_0_jtag_debug_module_readdata_from_sa                           (cpu_0_jtag_debug_module_readdata_from_sa),
      .d1_cpu_0_jtag_debug_module_end_xfer                                (d1_cpu_0_jtag_debug_module_end_xfer),
      .d1_nios_system_clock_2_in_end_xfer                                 (d1_nios_system_clock_2_in_end_xfer),
      .d1_onchip_memory2_0_s1_end_xfer                                    (d1_onchip_memory2_0_s1_end_xfer),
      .d1_onchip_memory2_1_s1_end_xfer                                    (d1_onchip_memory2_1_s1_end_xfer),
      .d1_onchip_memory2_2_s1_end_xfer                                    (d1_onchip_memory2_2_s1_end_xfer),
      .d1_onchip_memory2_3_s1_end_xfer                                    (d1_onchip_memory2_3_s1_end_xfer),
      .nios_system_clock_2_in_readdata_from_sa                            (nios_system_clock_2_in_readdata_from_sa),
      .nios_system_clock_2_in_waitrequest_from_sa                         (nios_system_clock_2_in_waitrequest_from_sa),
      .onchip_memory2_0_s1_readdata_from_sa                               (onchip_memory2_0_s1_readdata_from_sa),
      .onchip_memory2_1_s1_readdata_from_sa                               (onchip_memory2_1_s1_readdata_from_sa),
      .onchip_memory2_2_s1_readdata_from_sa                               (onchip_memory2_2_s1_readdata_from_sa),
      .onchip_memory2_3_s1_readdata_from_sa                               (onchip_memory2_3_s1_readdata_from_sa),
      .reset_n                                                            (sys_clk_reset_n)
    );

  cpu_0 the_cpu_0
    (
      .A_ci_multi_a                          (cpu_0_custom_instruction_master_multi_a),
      .A_ci_multi_b                          (cpu_0_custom_instruction_master_multi_b),
      .A_ci_multi_c                          (cpu_0_custom_instruction_master_multi_c),
      .A_ci_multi_clk_en                     (cpu_0_custom_instruction_master_multi_clk_en),
      .A_ci_multi_clock                      (cpu_0_custom_instruction_master_multi_clk),
      .A_ci_multi_dataa                      (cpu_0_custom_instruction_master_multi_dataa),
      .A_ci_multi_datab                      (cpu_0_custom_instruction_master_multi_datab),
      .A_ci_multi_done                       (cpu_0_custom_instruction_master_multi_done),
      .A_ci_multi_estatus                    (cpu_0_custom_instruction_master_multi_estatus),
      .A_ci_multi_ipending                   (cpu_0_custom_instruction_master_multi_ipending),
      .A_ci_multi_n                          (cpu_0_custom_instruction_master_multi_n),
      .A_ci_multi_readra                     (cpu_0_custom_instruction_master_multi_readra),
      .A_ci_multi_readrb                     (cpu_0_custom_instruction_master_multi_readrb),
      .A_ci_multi_reset                      (cpu_0_custom_instruction_master_multi_reset),
      .A_ci_multi_result                     (cpu_0_custom_instruction_master_multi_result),
      .A_ci_multi_start                      (cpu_0_custom_instruction_master_multi_start),
      .A_ci_multi_status                     (cpu_0_custom_instruction_master_multi_status),
      .A_ci_multi_writerc                    (cpu_0_custom_instruction_master_multi_writerc),
      .clk                                   (sys_clk),
      .d_address                             (cpu_0_data_master_address),
      .d_byteenable                          (cpu_0_data_master_byteenable),
      .d_irq                                 (cpu_0_data_master_irq),
      .d_read                                (cpu_0_data_master_read),
      .d_readdata                            (cpu_0_data_master_readdata),
      .d_readdatavalid                       (cpu_0_data_master_readdatavalid),
      .d_waitrequest                         (cpu_0_data_master_waitrequest),
      .d_write                               (cpu_0_data_master_write),
      .d_writedata                           (cpu_0_data_master_writedata),
      .i_address                             (cpu_0_instruction_master_address),
      .i_read                                (cpu_0_instruction_master_read),
      .i_readdata                            (cpu_0_instruction_master_readdata),
      .i_readdatavalid                       (cpu_0_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_0_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_0_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_0_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_0_jtag_debug_module_byteenable),
      .jtag_debug_module_debugaccess         (cpu_0_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_0_jtag_debug_module_readdata),
      .jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_0_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_0_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_0_jtag_debug_module_writedata),
      .reset_n                               (cpu_0_custom_instruction_master_reset_n)
    );

  cpu_0_altera_nios_custom_instr_floating_point_inst_s1_arbitrator the_cpu_0_altera_nios_custom_instr_floating_point_inst_s1
    (
      .clk                                                                                         (sys_clk),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_clk_en                                (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_clk_en),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_dataa                                 (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_dataa),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_datab                                 (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_datab),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done                                  (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa                          (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_n                                     (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_n),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_reset                                 (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_reset),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result                                (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa                        (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select                                (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_select),
      .cpu_0_altera_nios_custom_instr_floating_point_inst_s1_start                                 (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_start),
      .cpu_0_custom_instruction_master_multi_clk_en                                                (cpu_0_custom_instruction_master_multi_clk_en),
      .cpu_0_custom_instruction_master_multi_dataa                                                 (cpu_0_custom_instruction_master_multi_dataa),
      .cpu_0_custom_instruction_master_multi_datab                                                 (cpu_0_custom_instruction_master_multi_datab),
      .cpu_0_custom_instruction_master_multi_n                                                     (cpu_0_custom_instruction_master_multi_n),
      .cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1 (cpu_0_custom_instruction_master_start_cpu_0_altera_nios_custom_instr_floating_point_inst_s1),
      .reset_n                                                                                     (sys_clk_reset_n)
    );

  cpu_0_altera_nios_custom_instr_floating_point_inst the_cpu_0_altera_nios_custom_instr_floating_point_inst
    (
      .clk    (sys_clk),
      .clk_en (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_clk_en),
      .dataa  (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_dataa),
      .datab  (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_datab),
      .done   (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_done),
      .n      (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_n),
      .reset  (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_reset),
      .result (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_result),
      .start  (cpu_0_altera_nios_custom_instr_floating_point_inst_s1_start)
    );

  cpu_1_jtag_debug_module_arbitrator the_cpu_1_jtag_debug_module
    (
      .clk                                                                              (sys_clk),
      .cpu_1_data_master_address_to_slave                                               (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_byteenable                                                     (cpu_1_data_master_byteenable),
      .cpu_1_data_master_debugaccess                                                    (cpu_1_data_master_debugaccess),
      .cpu_1_data_master_granted_cpu_1_jtag_debug_module                                (cpu_1_data_master_granted_cpu_1_jtag_debug_module),
      .cpu_1_data_master_latency_counter                                                (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module                      (cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module),
      .cpu_1_data_master_read                                                           (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module                        (cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_cpu_1_jtag_debug_module                               (cpu_1_data_master_requests_cpu_1_jtag_debug_module),
      .cpu_1_data_master_write                                                          (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                                      (cpu_1_data_master_writedata),
      .cpu_1_instruction_master_address_to_slave                                        (cpu_1_instruction_master_address_to_slave),
      .cpu_1_instruction_master_granted_cpu_1_jtag_debug_module                         (cpu_1_instruction_master_granted_cpu_1_jtag_debug_module),
      .cpu_1_instruction_master_latency_counter                                         (cpu_1_instruction_master_latency_counter),
      .cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module               (cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module),
      .cpu_1_instruction_master_read                                                    (cpu_1_instruction_master_read),
      .cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module                 (cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module),
      .cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_instruction_master_requests_cpu_1_jtag_debug_module                        (cpu_1_instruction_master_requests_cpu_1_jtag_debug_module),
      .cpu_1_jtag_debug_module_address                                                  (cpu_1_jtag_debug_module_address),
      .cpu_1_jtag_debug_module_begintransfer                                            (cpu_1_jtag_debug_module_begintransfer),
      .cpu_1_jtag_debug_module_byteenable                                               (cpu_1_jtag_debug_module_byteenable),
      .cpu_1_jtag_debug_module_chipselect                                               (cpu_1_jtag_debug_module_chipselect),
      .cpu_1_jtag_debug_module_debugaccess                                              (cpu_1_jtag_debug_module_debugaccess),
      .cpu_1_jtag_debug_module_readdata                                                 (cpu_1_jtag_debug_module_readdata),
      .cpu_1_jtag_debug_module_readdata_from_sa                                         (cpu_1_jtag_debug_module_readdata_from_sa),
      .cpu_1_jtag_debug_module_resetrequest                                             (cpu_1_jtag_debug_module_resetrequest),
      .cpu_1_jtag_debug_module_resetrequest_from_sa                                     (cpu_1_jtag_debug_module_resetrequest_from_sa),
      .cpu_1_jtag_debug_module_write                                                    (cpu_1_jtag_debug_module_write),
      .cpu_1_jtag_debug_module_writedata                                                (cpu_1_jtag_debug_module_writedata),
      .d1_cpu_1_jtag_debug_module_end_xfer                                              (d1_cpu_1_jtag_debug_module_end_xfer),
      .reset_n                                                                          (sys_clk_reset_n)
    );

  cpu_1_custom_instruction_master_arbitrator the_cpu_1_custom_instruction_master
    (
      .clk                                                                                         (sys_clk),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa                          (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa                        (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select                                (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select),
      .cpu_1_custom_instruction_master_multi_done                                                  (cpu_1_custom_instruction_master_multi_done),
      .cpu_1_custom_instruction_master_multi_result                                                (cpu_1_custom_instruction_master_multi_result),
      .cpu_1_custom_instruction_master_multi_start                                                 (cpu_1_custom_instruction_master_multi_start),
      .cpu_1_custom_instruction_master_reset_n                                                     (cpu_1_custom_instruction_master_reset_n),
      .cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1 (cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1),
      .reset_n                                                                                     (sys_clk_reset_n)
    );

  cpu_1_data_master_arbitrator the_cpu_1_data_master
    (
      .clk                                                                               (sys_clk),
      .cpu_1_data_master_address                                                         (cpu_1_data_master_address),
      .cpu_1_data_master_address_to_slave                                                (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_byteenable                                                      (cpu_1_data_master_byteenable),
      .cpu_1_data_master_byteenable_nios_system_clock_1_in                               (cpu_1_data_master_byteenable_nios_system_clock_1_in),
      .cpu_1_data_master_byteenable_nios_system_clock_8_in                               (cpu_1_data_master_byteenable_nios_system_clock_8_in),
      .cpu_1_data_master_byteenable_sram_0_avalon_sram_slave                             (cpu_1_data_master_byteenable_sram_0_avalon_sram_slave),
      .cpu_1_data_master_dbs_address                                                     (cpu_1_data_master_dbs_address),
      .cpu_1_data_master_dbs_write_16                                                    (cpu_1_data_master_dbs_write_16),
      .cpu_1_data_master_dbs_write_8                                                     (cpu_1_data_master_dbs_write_8),
      .cpu_1_data_master_granted_cpu_1_jtag_debug_module                                 (cpu_1_data_master_granted_cpu_1_jtag_debug_module),
      .cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave                           (cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave),
      .cpu_1_data_master_granted_keys_s1                                                 (cpu_1_data_master_granted_keys_s1),
      .cpu_1_data_master_granted_mailbox_0_s1                                            (cpu_1_data_master_granted_mailbox_0_s1),
      .cpu_1_data_master_granted_mailbox_1_s1                                            (cpu_1_data_master_granted_mailbox_1_s1),
      .cpu_1_data_master_granted_mailbox_2_s1                                            (cpu_1_data_master_granted_mailbox_2_s1),
      .cpu_1_data_master_granted_mailbox_3_s1                                            (cpu_1_data_master_granted_mailbox_3_s1),
      .cpu_1_data_master_granted_nios_system_clock_1_in                                  (cpu_1_data_master_granted_nios_system_clock_1_in),
      .cpu_1_data_master_granted_nios_system_clock_8_in                                  (cpu_1_data_master_granted_nios_system_clock_8_in),
      .cpu_1_data_master_granted_onchip_memory2_0_s1                                     (cpu_1_data_master_granted_onchip_memory2_0_s1),
      .cpu_1_data_master_granted_onchip_memory2_1_s1                                     (cpu_1_data_master_granted_onchip_memory2_1_s1),
      .cpu_1_data_master_granted_onchip_memory2_2_s1                                     (cpu_1_data_master_granted_onchip_memory2_2_s1),
      .cpu_1_data_master_granted_onchip_memory2_3_s1                                     (cpu_1_data_master_granted_onchip_memory2_3_s1),
      .cpu_1_data_master_granted_performance_counter_0_control_slave                     (cpu_1_data_master_granted_performance_counter_0_control_slave),
      .cpu_1_data_master_granted_sram_0_avalon_sram_slave                                (cpu_1_data_master_granted_sram_0_avalon_sram_slave),
      .cpu_1_data_master_granted_sysid_control_slave                                     (cpu_1_data_master_granted_sysid_control_slave),
      .cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave           (cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_1_data_master_irq                                                             (cpu_1_data_master_irq),
      .cpu_1_data_master_latency_counter                                                 (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module                       (cpu_1_data_master_qualified_request_cpu_1_jtag_debug_module),
      .cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave                 (cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave),
      .cpu_1_data_master_qualified_request_keys_s1                                       (cpu_1_data_master_qualified_request_keys_s1),
      .cpu_1_data_master_qualified_request_mailbox_0_s1                                  (cpu_1_data_master_qualified_request_mailbox_0_s1),
      .cpu_1_data_master_qualified_request_mailbox_1_s1                                  (cpu_1_data_master_qualified_request_mailbox_1_s1),
      .cpu_1_data_master_qualified_request_mailbox_2_s1                                  (cpu_1_data_master_qualified_request_mailbox_2_s1),
      .cpu_1_data_master_qualified_request_mailbox_3_s1                                  (cpu_1_data_master_qualified_request_mailbox_3_s1),
      .cpu_1_data_master_qualified_request_nios_system_clock_1_in                        (cpu_1_data_master_qualified_request_nios_system_clock_1_in),
      .cpu_1_data_master_qualified_request_nios_system_clock_8_in                        (cpu_1_data_master_qualified_request_nios_system_clock_8_in),
      .cpu_1_data_master_qualified_request_onchip_memory2_0_s1                           (cpu_1_data_master_qualified_request_onchip_memory2_0_s1),
      .cpu_1_data_master_qualified_request_onchip_memory2_1_s1                           (cpu_1_data_master_qualified_request_onchip_memory2_1_s1),
      .cpu_1_data_master_qualified_request_onchip_memory2_2_s1                           (cpu_1_data_master_qualified_request_onchip_memory2_2_s1),
      .cpu_1_data_master_qualified_request_onchip_memory2_3_s1                           (cpu_1_data_master_qualified_request_onchip_memory2_3_s1),
      .cpu_1_data_master_qualified_request_performance_counter_0_control_slave           (cpu_1_data_master_qualified_request_performance_counter_0_control_slave),
      .cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave                      (cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_1_data_master_qualified_request_sysid_control_slave                           (cpu_1_data_master_qualified_request_sysid_control_slave),
      .cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave (cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_1_data_master_read                                                            (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module                         (cpu_1_data_master_read_data_valid_cpu_1_jtag_debug_module),
      .cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave                   (cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave),
      .cpu_1_data_master_read_data_valid_keys_s1                                         (cpu_1_data_master_read_data_valid_keys_s1),
      .cpu_1_data_master_read_data_valid_mailbox_0_s1                                    (cpu_1_data_master_read_data_valid_mailbox_0_s1),
      .cpu_1_data_master_read_data_valid_mailbox_1_s1                                    (cpu_1_data_master_read_data_valid_mailbox_1_s1),
      .cpu_1_data_master_read_data_valid_mailbox_2_s1                                    (cpu_1_data_master_read_data_valid_mailbox_2_s1),
      .cpu_1_data_master_read_data_valid_mailbox_3_s1                                    (cpu_1_data_master_read_data_valid_mailbox_3_s1),
      .cpu_1_data_master_read_data_valid_nios_system_clock_1_in                          (cpu_1_data_master_read_data_valid_nios_system_clock_1_in),
      .cpu_1_data_master_read_data_valid_nios_system_clock_8_in                          (cpu_1_data_master_read_data_valid_nios_system_clock_8_in),
      .cpu_1_data_master_read_data_valid_onchip_memory2_0_s1                             (cpu_1_data_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_1_data_master_read_data_valid_onchip_memory2_1_s1                             (cpu_1_data_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_1_data_master_read_data_valid_onchip_memory2_2_s1                             (cpu_1_data_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_1_data_master_read_data_valid_onchip_memory2_3_s1                             (cpu_1_data_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_1_data_master_read_data_valid_performance_counter_0_control_slave             (cpu_1_data_master_read_data_valid_performance_counter_0_control_slave),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave                        (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register         (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_read_data_valid_sysid_control_slave                             (cpu_1_data_master_read_data_valid_sysid_control_slave),
      .cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave   (cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_1_data_master_readdata                                                        (cpu_1_data_master_readdata),
      .cpu_1_data_master_readdatavalid                                                   (cpu_1_data_master_readdatavalid),
      .cpu_1_data_master_requests_cpu_1_jtag_debug_module                                (cpu_1_data_master_requests_cpu_1_jtag_debug_module),
      .cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave                          (cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave),
      .cpu_1_data_master_requests_keys_s1                                                (cpu_1_data_master_requests_keys_s1),
      .cpu_1_data_master_requests_mailbox_0_s1                                           (cpu_1_data_master_requests_mailbox_0_s1),
      .cpu_1_data_master_requests_mailbox_1_s1                                           (cpu_1_data_master_requests_mailbox_1_s1),
      .cpu_1_data_master_requests_mailbox_2_s1                                           (cpu_1_data_master_requests_mailbox_2_s1),
      .cpu_1_data_master_requests_mailbox_3_s1                                           (cpu_1_data_master_requests_mailbox_3_s1),
      .cpu_1_data_master_requests_nios_system_clock_1_in                                 (cpu_1_data_master_requests_nios_system_clock_1_in),
      .cpu_1_data_master_requests_nios_system_clock_8_in                                 (cpu_1_data_master_requests_nios_system_clock_8_in),
      .cpu_1_data_master_requests_onchip_memory2_0_s1                                    (cpu_1_data_master_requests_onchip_memory2_0_s1),
      .cpu_1_data_master_requests_onchip_memory2_1_s1                                    (cpu_1_data_master_requests_onchip_memory2_1_s1),
      .cpu_1_data_master_requests_onchip_memory2_2_s1                                    (cpu_1_data_master_requests_onchip_memory2_2_s1),
      .cpu_1_data_master_requests_onchip_memory2_3_s1                                    (cpu_1_data_master_requests_onchip_memory2_3_s1),
      .cpu_1_data_master_requests_performance_counter_0_control_slave                    (cpu_1_data_master_requests_performance_counter_0_control_slave),
      .cpu_1_data_master_requests_sram_0_avalon_sram_slave                               (cpu_1_data_master_requests_sram_0_avalon_sram_slave),
      .cpu_1_data_master_requests_sysid_control_slave                                    (cpu_1_data_master_requests_sysid_control_slave),
      .cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave          (cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_1_data_master_waitrequest                                                     (cpu_1_data_master_waitrequest),
      .cpu_1_data_master_write                                                           (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                                       (cpu_1_data_master_writedata),
      .cpu_1_jtag_debug_module_readdata_from_sa                                          (cpu_1_jtag_debug_module_readdata_from_sa),
      .d1_cpu_1_jtag_debug_module_end_xfer                                               (d1_cpu_1_jtag_debug_module_end_xfer),
      .d1_jtag_uart_1_avalon_jtag_slave_end_xfer                                         (d1_jtag_uart_1_avalon_jtag_slave_end_xfer),
      .d1_keys_s1_end_xfer                                                               (d1_keys_s1_end_xfer),
      .d1_mailbox_0_s1_end_xfer                                                          (d1_mailbox_0_s1_end_xfer),
      .d1_mailbox_1_s1_end_xfer                                                          (d1_mailbox_1_s1_end_xfer),
      .d1_mailbox_2_s1_end_xfer                                                          (d1_mailbox_2_s1_end_xfer),
      .d1_mailbox_3_s1_end_xfer                                                          (d1_mailbox_3_s1_end_xfer),
      .d1_nios_system_clock_1_in_end_xfer                                                (d1_nios_system_clock_1_in_end_xfer),
      .d1_nios_system_clock_8_in_end_xfer                                                (d1_nios_system_clock_8_in_end_xfer),
      .d1_onchip_memory2_0_s1_end_xfer                                                   (d1_onchip_memory2_0_s1_end_xfer),
      .d1_onchip_memory2_1_s1_end_xfer                                                   (d1_onchip_memory2_1_s1_end_xfer),
      .d1_onchip_memory2_2_s1_end_xfer                                                   (d1_onchip_memory2_2_s1_end_xfer),
      .d1_onchip_memory2_3_s1_end_xfer                                                   (d1_onchip_memory2_3_s1_end_xfer),
      .d1_performance_counter_0_control_slave_end_xfer                                   (d1_performance_counter_0_control_slave_end_xfer),
      .d1_sram_0_avalon_sram_slave_end_xfer                                              (d1_sram_0_avalon_sram_slave_end_xfer),
      .d1_sysid_control_slave_end_xfer                                                   (d1_sysid_control_slave_end_xfer),
      .d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer                         (d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer),
      .jtag_uart_1_avalon_jtag_slave_irq_from_sa                                         (jtag_uart_1_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_1_avalon_jtag_slave_readdata_from_sa                                    (jtag_uart_1_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa                                 (jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa),
      .keys_s1_readdata_from_sa                                                          (keys_s1_readdata_from_sa),
      .mailbox_0_s1_readdata_from_sa                                                     (mailbox_0_s1_readdata_from_sa),
      .mailbox_1_s1_readdata_from_sa                                                     (mailbox_1_s1_readdata_from_sa),
      .mailbox_2_s1_readdata_from_sa                                                     (mailbox_2_s1_readdata_from_sa),
      .mailbox_3_s1_readdata_from_sa                                                     (mailbox_3_s1_readdata_from_sa),
      .nios_system_clock_1_in_readdata_from_sa                                           (nios_system_clock_1_in_readdata_from_sa),
      .nios_system_clock_1_in_waitrequest_from_sa                                        (nios_system_clock_1_in_waitrequest_from_sa),
      .nios_system_clock_8_in_readdata_from_sa                                           (nios_system_clock_8_in_readdata_from_sa),
      .nios_system_clock_8_in_waitrequest_from_sa                                        (nios_system_clock_8_in_waitrequest_from_sa),
      .onchip_memory2_0_s1_readdata_from_sa                                              (onchip_memory2_0_s1_readdata_from_sa),
      .onchip_memory2_1_s1_readdata_from_sa                                              (onchip_memory2_1_s1_readdata_from_sa),
      .onchip_memory2_2_s1_readdata_from_sa                                              (onchip_memory2_2_s1_readdata_from_sa),
      .onchip_memory2_3_s1_readdata_from_sa                                              (onchip_memory2_3_s1_readdata_from_sa),
      .performance_counter_0_control_slave_readdata_from_sa                              (performance_counter_0_control_slave_readdata_from_sa),
      .reset_n                                                                           (sys_clk_reset_n),
      .sram_0_avalon_sram_slave_readdata_from_sa                                         (sram_0_avalon_sram_slave_readdata_from_sa),
      .sysid_control_slave_readdata_from_sa                                              (sysid_control_slave_readdata_from_sa),
      .video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa                    (video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa)
    );

  cpu_1_instruction_master_arbitrator the_cpu_1_instruction_master
    (
      .clk                                                                              (sys_clk),
      .cpu_1_instruction_master_address                                                 (cpu_1_instruction_master_address),
      .cpu_1_instruction_master_address_to_slave                                        (cpu_1_instruction_master_address_to_slave),
      .cpu_1_instruction_master_dbs_address                                             (cpu_1_instruction_master_dbs_address),
      .cpu_1_instruction_master_granted_cpu_1_jtag_debug_module                         (cpu_1_instruction_master_granted_cpu_1_jtag_debug_module),
      .cpu_1_instruction_master_granted_nios_system_clock_0_in                          (cpu_1_instruction_master_granted_nios_system_clock_0_in),
      .cpu_1_instruction_master_granted_onchip_memory2_0_s1                             (cpu_1_instruction_master_granted_onchip_memory2_0_s1),
      .cpu_1_instruction_master_granted_onchip_memory2_1_s1                             (cpu_1_instruction_master_granted_onchip_memory2_1_s1),
      .cpu_1_instruction_master_granted_onchip_memory2_2_s1                             (cpu_1_instruction_master_granted_onchip_memory2_2_s1),
      .cpu_1_instruction_master_granted_onchip_memory2_3_s1                             (cpu_1_instruction_master_granted_onchip_memory2_3_s1),
      .cpu_1_instruction_master_granted_sram_0_avalon_sram_slave                        (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave),
      .cpu_1_instruction_master_latency_counter                                         (cpu_1_instruction_master_latency_counter),
      .cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module               (cpu_1_instruction_master_qualified_request_cpu_1_jtag_debug_module),
      .cpu_1_instruction_master_qualified_request_nios_system_clock_0_in                (cpu_1_instruction_master_qualified_request_nios_system_clock_0_in),
      .cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1                   (cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1),
      .cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1                   (cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1),
      .cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1                   (cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1),
      .cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1                   (cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1),
      .cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave              (cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_1_instruction_master_read                                                    (cpu_1_instruction_master_read),
      .cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module                 (cpu_1_instruction_master_read_data_valid_cpu_1_jtag_debug_module),
      .cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in                  (cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in),
      .cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1                     (cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1                     (cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1                     (cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1                     (cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave                (cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_instruction_master_readdata                                                (cpu_1_instruction_master_readdata),
      .cpu_1_instruction_master_readdatavalid                                           (cpu_1_instruction_master_readdatavalid),
      .cpu_1_instruction_master_requests_cpu_1_jtag_debug_module                        (cpu_1_instruction_master_requests_cpu_1_jtag_debug_module),
      .cpu_1_instruction_master_requests_nios_system_clock_0_in                         (cpu_1_instruction_master_requests_nios_system_clock_0_in),
      .cpu_1_instruction_master_requests_onchip_memory2_0_s1                            (cpu_1_instruction_master_requests_onchip_memory2_0_s1),
      .cpu_1_instruction_master_requests_onchip_memory2_1_s1                            (cpu_1_instruction_master_requests_onchip_memory2_1_s1),
      .cpu_1_instruction_master_requests_onchip_memory2_2_s1                            (cpu_1_instruction_master_requests_onchip_memory2_2_s1),
      .cpu_1_instruction_master_requests_onchip_memory2_3_s1                            (cpu_1_instruction_master_requests_onchip_memory2_3_s1),
      .cpu_1_instruction_master_requests_sram_0_avalon_sram_slave                       (cpu_1_instruction_master_requests_sram_0_avalon_sram_slave),
      .cpu_1_instruction_master_waitrequest                                             (cpu_1_instruction_master_waitrequest),
      .cpu_1_jtag_debug_module_readdata_from_sa                                         (cpu_1_jtag_debug_module_readdata_from_sa),
      .d1_cpu_1_jtag_debug_module_end_xfer                                              (d1_cpu_1_jtag_debug_module_end_xfer),
      .d1_nios_system_clock_0_in_end_xfer                                               (d1_nios_system_clock_0_in_end_xfer),
      .d1_onchip_memory2_0_s1_end_xfer                                                  (d1_onchip_memory2_0_s1_end_xfer),
      .d1_onchip_memory2_1_s1_end_xfer                                                  (d1_onchip_memory2_1_s1_end_xfer),
      .d1_onchip_memory2_2_s1_end_xfer                                                  (d1_onchip_memory2_2_s1_end_xfer),
      .d1_onchip_memory2_3_s1_end_xfer                                                  (d1_onchip_memory2_3_s1_end_xfer),
      .d1_sram_0_avalon_sram_slave_end_xfer                                             (d1_sram_0_avalon_sram_slave_end_xfer),
      .nios_system_clock_0_in_readdata_from_sa                                          (nios_system_clock_0_in_readdata_from_sa),
      .nios_system_clock_0_in_waitrequest_from_sa                                       (nios_system_clock_0_in_waitrequest_from_sa),
      .onchip_memory2_0_s1_readdata_from_sa                                             (onchip_memory2_0_s1_readdata_from_sa),
      .onchip_memory2_1_s1_readdata_from_sa                                             (onchip_memory2_1_s1_readdata_from_sa),
      .onchip_memory2_2_s1_readdata_from_sa                                             (onchip_memory2_2_s1_readdata_from_sa),
      .onchip_memory2_3_s1_readdata_from_sa                                             (onchip_memory2_3_s1_readdata_from_sa),
      .reset_n                                                                          (sys_clk_reset_n),
      .sram_0_avalon_sram_slave_readdata_from_sa                                        (sram_0_avalon_sram_slave_readdata_from_sa)
    );

  cpu_1 the_cpu_1
    (
      .A_ci_multi_a                          (cpu_1_custom_instruction_master_multi_a),
      .A_ci_multi_b                          (cpu_1_custom_instruction_master_multi_b),
      .A_ci_multi_c                          (cpu_1_custom_instruction_master_multi_c),
      .A_ci_multi_clk_en                     (cpu_1_custom_instruction_master_multi_clk_en),
      .A_ci_multi_clock                      (cpu_1_custom_instruction_master_multi_clk),
      .A_ci_multi_dataa                      (cpu_1_custom_instruction_master_multi_dataa),
      .A_ci_multi_datab                      (cpu_1_custom_instruction_master_multi_datab),
      .A_ci_multi_done                       (cpu_1_custom_instruction_master_multi_done),
      .A_ci_multi_estatus                    (cpu_1_custom_instruction_master_multi_estatus),
      .A_ci_multi_ipending                   (cpu_1_custom_instruction_master_multi_ipending),
      .A_ci_multi_n                          (cpu_1_custom_instruction_master_multi_n),
      .A_ci_multi_readra                     (cpu_1_custom_instruction_master_multi_readra),
      .A_ci_multi_readrb                     (cpu_1_custom_instruction_master_multi_readrb),
      .A_ci_multi_reset                      (cpu_1_custom_instruction_master_multi_reset),
      .A_ci_multi_result                     (cpu_1_custom_instruction_master_multi_result),
      .A_ci_multi_start                      (cpu_1_custom_instruction_master_multi_start),
      .A_ci_multi_status                     (cpu_1_custom_instruction_master_multi_status),
      .A_ci_multi_writerc                    (cpu_1_custom_instruction_master_multi_writerc),
      .clk                                   (sys_clk),
      .d_address                             (cpu_1_data_master_address),
      .d_byteenable                          (cpu_1_data_master_byteenable),
      .d_irq                                 (cpu_1_data_master_irq),
      .d_read                                (cpu_1_data_master_read),
      .d_readdata                            (cpu_1_data_master_readdata),
      .d_readdatavalid                       (cpu_1_data_master_readdatavalid),
      .d_waitrequest                         (cpu_1_data_master_waitrequest),
      .d_write                               (cpu_1_data_master_write),
      .d_writedata                           (cpu_1_data_master_writedata),
      .i_address                             (cpu_1_instruction_master_address),
      .i_read                                (cpu_1_instruction_master_read),
      .i_readdata                            (cpu_1_instruction_master_readdata),
      .i_readdatavalid                       (cpu_1_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_1_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_1_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_1_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_1_jtag_debug_module_byteenable),
      .jtag_debug_module_debugaccess         (cpu_1_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_1_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_1_jtag_debug_module_readdata),
      .jtag_debug_module_resetrequest        (cpu_1_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_1_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_1_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_1_jtag_debug_module_writedata),
      .reset_n                               (cpu_1_custom_instruction_master_reset_n)
    );

  cpu_1_altera_nios_custom_instr_floating_point_inst_s1_arbitrator the_cpu_1_altera_nios_custom_instr_floating_point_inst_s1
    (
      .clk                                                                                         (sys_clk),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_clk_en                                (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_clk_en),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_dataa                                 (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_dataa),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_datab                                 (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_datab),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done                                  (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa                          (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_n                                     (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_n),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_reset                                 (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_reset),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result                                (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa                        (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select                                (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_select),
      .cpu_1_altera_nios_custom_instr_floating_point_inst_s1_start                                 (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_start),
      .cpu_1_custom_instruction_master_multi_clk_en                                                (cpu_1_custom_instruction_master_multi_clk_en),
      .cpu_1_custom_instruction_master_multi_dataa                                                 (cpu_1_custom_instruction_master_multi_dataa),
      .cpu_1_custom_instruction_master_multi_datab                                                 (cpu_1_custom_instruction_master_multi_datab),
      .cpu_1_custom_instruction_master_multi_n                                                     (cpu_1_custom_instruction_master_multi_n),
      .cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1 (cpu_1_custom_instruction_master_start_cpu_1_altera_nios_custom_instr_floating_point_inst_s1),
      .reset_n                                                                                     (sys_clk_reset_n)
    );

  cpu_1_altera_nios_custom_instr_floating_point_inst the_cpu_1_altera_nios_custom_instr_floating_point_inst
    (
      .clk    (sys_clk),
      .clk_en (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_clk_en),
      .dataa  (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_dataa),
      .datab  (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_datab),
      .done   (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_done),
      .n      (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_n),
      .reset  (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_reset),
      .result (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_result),
      .start  (cpu_1_altera_nios_custom_instr_floating_point_inst_s1_start)
    );

  cpu_2_jtag_debug_module_arbitrator the_cpu_2_jtag_debug_module
    (
      .clk                                                                              (sys_clk),
      .cpu_2_data_master_address_to_slave                                               (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_byteenable                                                     (cpu_2_data_master_byteenable),
      .cpu_2_data_master_debugaccess                                                    (cpu_2_data_master_debugaccess),
      .cpu_2_data_master_granted_cpu_2_jtag_debug_module                                (cpu_2_data_master_granted_cpu_2_jtag_debug_module),
      .cpu_2_data_master_latency_counter                                                (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module                      (cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module),
      .cpu_2_data_master_read                                                           (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module                        (cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_cpu_2_jtag_debug_module                               (cpu_2_data_master_requests_cpu_2_jtag_debug_module),
      .cpu_2_data_master_write                                                          (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                                      (cpu_2_data_master_writedata),
      .cpu_2_instruction_master_address_to_slave                                        (cpu_2_instruction_master_address_to_slave),
      .cpu_2_instruction_master_granted_cpu_2_jtag_debug_module                         (cpu_2_instruction_master_granted_cpu_2_jtag_debug_module),
      .cpu_2_instruction_master_latency_counter                                         (cpu_2_instruction_master_latency_counter),
      .cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module               (cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module),
      .cpu_2_instruction_master_read                                                    (cpu_2_instruction_master_read),
      .cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module                 (cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module),
      .cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_instruction_master_requests_cpu_2_jtag_debug_module                        (cpu_2_instruction_master_requests_cpu_2_jtag_debug_module),
      .cpu_2_jtag_debug_module_address                                                  (cpu_2_jtag_debug_module_address),
      .cpu_2_jtag_debug_module_begintransfer                                            (cpu_2_jtag_debug_module_begintransfer),
      .cpu_2_jtag_debug_module_byteenable                                               (cpu_2_jtag_debug_module_byteenable),
      .cpu_2_jtag_debug_module_chipselect                                               (cpu_2_jtag_debug_module_chipselect),
      .cpu_2_jtag_debug_module_debugaccess                                              (cpu_2_jtag_debug_module_debugaccess),
      .cpu_2_jtag_debug_module_readdata                                                 (cpu_2_jtag_debug_module_readdata),
      .cpu_2_jtag_debug_module_readdata_from_sa                                         (cpu_2_jtag_debug_module_readdata_from_sa),
      .cpu_2_jtag_debug_module_resetrequest                                             (cpu_2_jtag_debug_module_resetrequest),
      .cpu_2_jtag_debug_module_resetrequest_from_sa                                     (cpu_2_jtag_debug_module_resetrequest_from_sa),
      .cpu_2_jtag_debug_module_write                                                    (cpu_2_jtag_debug_module_write),
      .cpu_2_jtag_debug_module_writedata                                                (cpu_2_jtag_debug_module_writedata),
      .d1_cpu_2_jtag_debug_module_end_xfer                                              (d1_cpu_2_jtag_debug_module_end_xfer),
      .reset_n                                                                          (sys_clk_reset_n)
    );

  cpu_2_custom_instruction_master_arbitrator the_cpu_2_custom_instruction_master
    (
      .clk                                                                                         (sys_clk),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa                          (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa                        (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select                                (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select),
      .cpu_2_custom_instruction_master_multi_done                                                  (cpu_2_custom_instruction_master_multi_done),
      .cpu_2_custom_instruction_master_multi_result                                                (cpu_2_custom_instruction_master_multi_result),
      .cpu_2_custom_instruction_master_multi_start                                                 (cpu_2_custom_instruction_master_multi_start),
      .cpu_2_custom_instruction_master_reset_n                                                     (cpu_2_custom_instruction_master_reset_n),
      .cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1 (cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1),
      .reset_n                                                                                     (sys_clk_reset_n)
    );

  cpu_2_data_master_arbitrator the_cpu_2_data_master
    (
      .clk                                                                               (sys_clk),
      .cpu_2_data_master_address                                                         (cpu_2_data_master_address),
      .cpu_2_data_master_address_to_slave                                                (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_byteenable                                                      (cpu_2_data_master_byteenable),
      .cpu_2_data_master_byteenable_nios_system_clock_10_in                              (cpu_2_data_master_byteenable_nios_system_clock_10_in),
      .cpu_2_data_master_byteenable_nios_system_clock_5_in                               (cpu_2_data_master_byteenable_nios_system_clock_5_in),
      .cpu_2_data_master_byteenable_sram_0_avalon_sram_slave                             (cpu_2_data_master_byteenable_sram_0_avalon_sram_slave),
      .cpu_2_data_master_dbs_address                                                     (cpu_2_data_master_dbs_address),
      .cpu_2_data_master_dbs_write_16                                                    (cpu_2_data_master_dbs_write_16),
      .cpu_2_data_master_dbs_write_8                                                     (cpu_2_data_master_dbs_write_8),
      .cpu_2_data_master_granted_cpu_2_jtag_debug_module                                 (cpu_2_data_master_granted_cpu_2_jtag_debug_module),
      .cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave                           (cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave),
      .cpu_2_data_master_granted_keys_s1                                                 (cpu_2_data_master_granted_keys_s1),
      .cpu_2_data_master_granted_mailbox_0_s1                                            (cpu_2_data_master_granted_mailbox_0_s1),
      .cpu_2_data_master_granted_mailbox_1_s1                                            (cpu_2_data_master_granted_mailbox_1_s1),
      .cpu_2_data_master_granted_mailbox_2_s1                                            (cpu_2_data_master_granted_mailbox_2_s1),
      .cpu_2_data_master_granted_mailbox_3_s1                                            (cpu_2_data_master_granted_mailbox_3_s1),
      .cpu_2_data_master_granted_nios_system_clock_10_in                                 (cpu_2_data_master_granted_nios_system_clock_10_in),
      .cpu_2_data_master_granted_nios_system_clock_5_in                                  (cpu_2_data_master_granted_nios_system_clock_5_in),
      .cpu_2_data_master_granted_onchip_memory2_0_s1                                     (cpu_2_data_master_granted_onchip_memory2_0_s1),
      .cpu_2_data_master_granted_onchip_memory2_1_s1                                     (cpu_2_data_master_granted_onchip_memory2_1_s1),
      .cpu_2_data_master_granted_onchip_memory2_2_s1                                     (cpu_2_data_master_granted_onchip_memory2_2_s1),
      .cpu_2_data_master_granted_onchip_memory2_3_s1                                     (cpu_2_data_master_granted_onchip_memory2_3_s1),
      .cpu_2_data_master_granted_performance_counter_0_control_slave                     (cpu_2_data_master_granted_performance_counter_0_control_slave),
      .cpu_2_data_master_granted_sram_0_avalon_sram_slave                                (cpu_2_data_master_granted_sram_0_avalon_sram_slave),
      .cpu_2_data_master_granted_sysid_control_slave                                     (cpu_2_data_master_granted_sysid_control_slave),
      .cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave           (cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_2_data_master_irq                                                             (cpu_2_data_master_irq),
      .cpu_2_data_master_latency_counter                                                 (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module                       (cpu_2_data_master_qualified_request_cpu_2_jtag_debug_module),
      .cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave                 (cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave),
      .cpu_2_data_master_qualified_request_keys_s1                                       (cpu_2_data_master_qualified_request_keys_s1),
      .cpu_2_data_master_qualified_request_mailbox_0_s1                                  (cpu_2_data_master_qualified_request_mailbox_0_s1),
      .cpu_2_data_master_qualified_request_mailbox_1_s1                                  (cpu_2_data_master_qualified_request_mailbox_1_s1),
      .cpu_2_data_master_qualified_request_mailbox_2_s1                                  (cpu_2_data_master_qualified_request_mailbox_2_s1),
      .cpu_2_data_master_qualified_request_mailbox_3_s1                                  (cpu_2_data_master_qualified_request_mailbox_3_s1),
      .cpu_2_data_master_qualified_request_nios_system_clock_10_in                       (cpu_2_data_master_qualified_request_nios_system_clock_10_in),
      .cpu_2_data_master_qualified_request_nios_system_clock_5_in                        (cpu_2_data_master_qualified_request_nios_system_clock_5_in),
      .cpu_2_data_master_qualified_request_onchip_memory2_0_s1                           (cpu_2_data_master_qualified_request_onchip_memory2_0_s1),
      .cpu_2_data_master_qualified_request_onchip_memory2_1_s1                           (cpu_2_data_master_qualified_request_onchip_memory2_1_s1),
      .cpu_2_data_master_qualified_request_onchip_memory2_2_s1                           (cpu_2_data_master_qualified_request_onchip_memory2_2_s1),
      .cpu_2_data_master_qualified_request_onchip_memory2_3_s1                           (cpu_2_data_master_qualified_request_onchip_memory2_3_s1),
      .cpu_2_data_master_qualified_request_performance_counter_0_control_slave           (cpu_2_data_master_qualified_request_performance_counter_0_control_slave),
      .cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave                      (cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_2_data_master_qualified_request_sysid_control_slave                           (cpu_2_data_master_qualified_request_sysid_control_slave),
      .cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave (cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_2_data_master_read                                                            (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module                         (cpu_2_data_master_read_data_valid_cpu_2_jtag_debug_module),
      .cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave                   (cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave),
      .cpu_2_data_master_read_data_valid_keys_s1                                         (cpu_2_data_master_read_data_valid_keys_s1),
      .cpu_2_data_master_read_data_valid_mailbox_0_s1                                    (cpu_2_data_master_read_data_valid_mailbox_0_s1),
      .cpu_2_data_master_read_data_valid_mailbox_1_s1                                    (cpu_2_data_master_read_data_valid_mailbox_1_s1),
      .cpu_2_data_master_read_data_valid_mailbox_2_s1                                    (cpu_2_data_master_read_data_valid_mailbox_2_s1),
      .cpu_2_data_master_read_data_valid_mailbox_3_s1                                    (cpu_2_data_master_read_data_valid_mailbox_3_s1),
      .cpu_2_data_master_read_data_valid_nios_system_clock_10_in                         (cpu_2_data_master_read_data_valid_nios_system_clock_10_in),
      .cpu_2_data_master_read_data_valid_nios_system_clock_5_in                          (cpu_2_data_master_read_data_valid_nios_system_clock_5_in),
      .cpu_2_data_master_read_data_valid_onchip_memory2_0_s1                             (cpu_2_data_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_2_data_master_read_data_valid_onchip_memory2_1_s1                             (cpu_2_data_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_2_data_master_read_data_valid_onchip_memory2_2_s1                             (cpu_2_data_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_2_data_master_read_data_valid_onchip_memory2_3_s1                             (cpu_2_data_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_2_data_master_read_data_valid_performance_counter_0_control_slave             (cpu_2_data_master_read_data_valid_performance_counter_0_control_slave),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave                        (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register         (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_read_data_valid_sysid_control_slave                             (cpu_2_data_master_read_data_valid_sysid_control_slave),
      .cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave   (cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_2_data_master_readdata                                                        (cpu_2_data_master_readdata),
      .cpu_2_data_master_readdatavalid                                                   (cpu_2_data_master_readdatavalid),
      .cpu_2_data_master_requests_cpu_2_jtag_debug_module                                (cpu_2_data_master_requests_cpu_2_jtag_debug_module),
      .cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave                          (cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave),
      .cpu_2_data_master_requests_keys_s1                                                (cpu_2_data_master_requests_keys_s1),
      .cpu_2_data_master_requests_mailbox_0_s1                                           (cpu_2_data_master_requests_mailbox_0_s1),
      .cpu_2_data_master_requests_mailbox_1_s1                                           (cpu_2_data_master_requests_mailbox_1_s1),
      .cpu_2_data_master_requests_mailbox_2_s1                                           (cpu_2_data_master_requests_mailbox_2_s1),
      .cpu_2_data_master_requests_mailbox_3_s1                                           (cpu_2_data_master_requests_mailbox_3_s1),
      .cpu_2_data_master_requests_nios_system_clock_10_in                                (cpu_2_data_master_requests_nios_system_clock_10_in),
      .cpu_2_data_master_requests_nios_system_clock_5_in                                 (cpu_2_data_master_requests_nios_system_clock_5_in),
      .cpu_2_data_master_requests_onchip_memory2_0_s1                                    (cpu_2_data_master_requests_onchip_memory2_0_s1),
      .cpu_2_data_master_requests_onchip_memory2_1_s1                                    (cpu_2_data_master_requests_onchip_memory2_1_s1),
      .cpu_2_data_master_requests_onchip_memory2_2_s1                                    (cpu_2_data_master_requests_onchip_memory2_2_s1),
      .cpu_2_data_master_requests_onchip_memory2_3_s1                                    (cpu_2_data_master_requests_onchip_memory2_3_s1),
      .cpu_2_data_master_requests_performance_counter_0_control_slave                    (cpu_2_data_master_requests_performance_counter_0_control_slave),
      .cpu_2_data_master_requests_sram_0_avalon_sram_slave                               (cpu_2_data_master_requests_sram_0_avalon_sram_slave),
      .cpu_2_data_master_requests_sysid_control_slave                                    (cpu_2_data_master_requests_sysid_control_slave),
      .cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave          (cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_2_data_master_waitrequest                                                     (cpu_2_data_master_waitrequest),
      .cpu_2_data_master_write                                                           (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                                       (cpu_2_data_master_writedata),
      .cpu_2_jtag_debug_module_readdata_from_sa                                          (cpu_2_jtag_debug_module_readdata_from_sa),
      .d1_cpu_2_jtag_debug_module_end_xfer                                               (d1_cpu_2_jtag_debug_module_end_xfer),
      .d1_jtag_uart_2_avalon_jtag_slave_end_xfer                                         (d1_jtag_uart_2_avalon_jtag_slave_end_xfer),
      .d1_keys_s1_end_xfer                                                               (d1_keys_s1_end_xfer),
      .d1_mailbox_0_s1_end_xfer                                                          (d1_mailbox_0_s1_end_xfer),
      .d1_mailbox_1_s1_end_xfer                                                          (d1_mailbox_1_s1_end_xfer),
      .d1_mailbox_2_s1_end_xfer                                                          (d1_mailbox_2_s1_end_xfer),
      .d1_mailbox_3_s1_end_xfer                                                          (d1_mailbox_3_s1_end_xfer),
      .d1_nios_system_clock_10_in_end_xfer                                               (d1_nios_system_clock_10_in_end_xfer),
      .d1_nios_system_clock_5_in_end_xfer                                                (d1_nios_system_clock_5_in_end_xfer),
      .d1_onchip_memory2_0_s1_end_xfer                                                   (d1_onchip_memory2_0_s1_end_xfer),
      .d1_onchip_memory2_1_s1_end_xfer                                                   (d1_onchip_memory2_1_s1_end_xfer),
      .d1_onchip_memory2_2_s1_end_xfer                                                   (d1_onchip_memory2_2_s1_end_xfer),
      .d1_onchip_memory2_3_s1_end_xfer                                                   (d1_onchip_memory2_3_s1_end_xfer),
      .d1_performance_counter_0_control_slave_end_xfer                                   (d1_performance_counter_0_control_slave_end_xfer),
      .d1_sram_0_avalon_sram_slave_end_xfer                                              (d1_sram_0_avalon_sram_slave_end_xfer),
      .d1_sysid_control_slave_end_xfer                                                   (d1_sysid_control_slave_end_xfer),
      .d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer                         (d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer),
      .jtag_uart_2_avalon_jtag_slave_irq_from_sa                                         (jtag_uart_2_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_2_avalon_jtag_slave_readdata_from_sa                                    (jtag_uart_2_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa                                 (jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa),
      .keys_s1_readdata_from_sa                                                          (keys_s1_readdata_from_sa),
      .mailbox_0_s1_readdata_from_sa                                                     (mailbox_0_s1_readdata_from_sa),
      .mailbox_1_s1_readdata_from_sa                                                     (mailbox_1_s1_readdata_from_sa),
      .mailbox_2_s1_readdata_from_sa                                                     (mailbox_2_s1_readdata_from_sa),
      .mailbox_3_s1_readdata_from_sa                                                     (mailbox_3_s1_readdata_from_sa),
      .nios_system_clock_10_in_readdata_from_sa                                          (nios_system_clock_10_in_readdata_from_sa),
      .nios_system_clock_10_in_waitrequest_from_sa                                       (nios_system_clock_10_in_waitrequest_from_sa),
      .nios_system_clock_5_in_readdata_from_sa                                           (nios_system_clock_5_in_readdata_from_sa),
      .nios_system_clock_5_in_waitrequest_from_sa                                        (nios_system_clock_5_in_waitrequest_from_sa),
      .onchip_memory2_0_s1_readdata_from_sa                                              (onchip_memory2_0_s1_readdata_from_sa),
      .onchip_memory2_1_s1_readdata_from_sa                                              (onchip_memory2_1_s1_readdata_from_sa),
      .onchip_memory2_2_s1_readdata_from_sa                                              (onchip_memory2_2_s1_readdata_from_sa),
      .onchip_memory2_3_s1_readdata_from_sa                                              (onchip_memory2_3_s1_readdata_from_sa),
      .performance_counter_0_control_slave_readdata_from_sa                              (performance_counter_0_control_slave_readdata_from_sa),
      .reset_n                                                                           (sys_clk_reset_n),
      .sram_0_avalon_sram_slave_readdata_from_sa                                         (sram_0_avalon_sram_slave_readdata_from_sa),
      .sysid_control_slave_readdata_from_sa                                              (sysid_control_slave_readdata_from_sa),
      .video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa                    (video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa)
    );

  cpu_2_instruction_master_arbitrator the_cpu_2_instruction_master
    (
      .clk                                                                              (sys_clk),
      .cpu_2_instruction_master_address                                                 (cpu_2_instruction_master_address),
      .cpu_2_instruction_master_address_to_slave                                        (cpu_2_instruction_master_address_to_slave),
      .cpu_2_instruction_master_dbs_address                                             (cpu_2_instruction_master_dbs_address),
      .cpu_2_instruction_master_granted_cpu_2_jtag_debug_module                         (cpu_2_instruction_master_granted_cpu_2_jtag_debug_module),
      .cpu_2_instruction_master_granted_nios_system_clock_4_in                          (cpu_2_instruction_master_granted_nios_system_clock_4_in),
      .cpu_2_instruction_master_granted_onchip_memory2_0_s1                             (cpu_2_instruction_master_granted_onchip_memory2_0_s1),
      .cpu_2_instruction_master_granted_onchip_memory2_1_s1                             (cpu_2_instruction_master_granted_onchip_memory2_1_s1),
      .cpu_2_instruction_master_granted_onchip_memory2_2_s1                             (cpu_2_instruction_master_granted_onchip_memory2_2_s1),
      .cpu_2_instruction_master_granted_onchip_memory2_3_s1                             (cpu_2_instruction_master_granted_onchip_memory2_3_s1),
      .cpu_2_instruction_master_granted_sram_0_avalon_sram_slave                        (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave),
      .cpu_2_instruction_master_latency_counter                                         (cpu_2_instruction_master_latency_counter),
      .cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module               (cpu_2_instruction_master_qualified_request_cpu_2_jtag_debug_module),
      .cpu_2_instruction_master_qualified_request_nios_system_clock_4_in                (cpu_2_instruction_master_qualified_request_nios_system_clock_4_in),
      .cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1                   (cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1),
      .cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1                   (cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1),
      .cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1                   (cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1),
      .cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1                   (cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1),
      .cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave              (cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_2_instruction_master_read                                                    (cpu_2_instruction_master_read),
      .cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module                 (cpu_2_instruction_master_read_data_valid_cpu_2_jtag_debug_module),
      .cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in                  (cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in),
      .cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1                     (cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1                     (cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1                     (cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1                     (cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave                (cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_instruction_master_readdata                                                (cpu_2_instruction_master_readdata),
      .cpu_2_instruction_master_readdatavalid                                           (cpu_2_instruction_master_readdatavalid),
      .cpu_2_instruction_master_requests_cpu_2_jtag_debug_module                        (cpu_2_instruction_master_requests_cpu_2_jtag_debug_module),
      .cpu_2_instruction_master_requests_nios_system_clock_4_in                         (cpu_2_instruction_master_requests_nios_system_clock_4_in),
      .cpu_2_instruction_master_requests_onchip_memory2_0_s1                            (cpu_2_instruction_master_requests_onchip_memory2_0_s1),
      .cpu_2_instruction_master_requests_onchip_memory2_1_s1                            (cpu_2_instruction_master_requests_onchip_memory2_1_s1),
      .cpu_2_instruction_master_requests_onchip_memory2_2_s1                            (cpu_2_instruction_master_requests_onchip_memory2_2_s1),
      .cpu_2_instruction_master_requests_onchip_memory2_3_s1                            (cpu_2_instruction_master_requests_onchip_memory2_3_s1),
      .cpu_2_instruction_master_requests_sram_0_avalon_sram_slave                       (cpu_2_instruction_master_requests_sram_0_avalon_sram_slave),
      .cpu_2_instruction_master_waitrequest                                             (cpu_2_instruction_master_waitrequest),
      .cpu_2_jtag_debug_module_readdata_from_sa                                         (cpu_2_jtag_debug_module_readdata_from_sa),
      .d1_cpu_2_jtag_debug_module_end_xfer                                              (d1_cpu_2_jtag_debug_module_end_xfer),
      .d1_nios_system_clock_4_in_end_xfer                                               (d1_nios_system_clock_4_in_end_xfer),
      .d1_onchip_memory2_0_s1_end_xfer                                                  (d1_onchip_memory2_0_s1_end_xfer),
      .d1_onchip_memory2_1_s1_end_xfer                                                  (d1_onchip_memory2_1_s1_end_xfer),
      .d1_onchip_memory2_2_s1_end_xfer                                                  (d1_onchip_memory2_2_s1_end_xfer),
      .d1_onchip_memory2_3_s1_end_xfer                                                  (d1_onchip_memory2_3_s1_end_xfer),
      .d1_sram_0_avalon_sram_slave_end_xfer                                             (d1_sram_0_avalon_sram_slave_end_xfer),
      .nios_system_clock_4_in_readdata_from_sa                                          (nios_system_clock_4_in_readdata_from_sa),
      .nios_system_clock_4_in_waitrequest_from_sa                                       (nios_system_clock_4_in_waitrequest_from_sa),
      .onchip_memory2_0_s1_readdata_from_sa                                             (onchip_memory2_0_s1_readdata_from_sa),
      .onchip_memory2_1_s1_readdata_from_sa                                             (onchip_memory2_1_s1_readdata_from_sa),
      .onchip_memory2_2_s1_readdata_from_sa                                             (onchip_memory2_2_s1_readdata_from_sa),
      .onchip_memory2_3_s1_readdata_from_sa                                             (onchip_memory2_3_s1_readdata_from_sa),
      .reset_n                                                                          (sys_clk_reset_n),
      .sram_0_avalon_sram_slave_readdata_from_sa                                        (sram_0_avalon_sram_slave_readdata_from_sa)
    );

  cpu_2 the_cpu_2
    (
      .A_ci_multi_a                          (cpu_2_custom_instruction_master_multi_a),
      .A_ci_multi_b                          (cpu_2_custom_instruction_master_multi_b),
      .A_ci_multi_c                          (cpu_2_custom_instruction_master_multi_c),
      .A_ci_multi_clk_en                     (cpu_2_custom_instruction_master_multi_clk_en),
      .A_ci_multi_clock                      (cpu_2_custom_instruction_master_multi_clk),
      .A_ci_multi_dataa                      (cpu_2_custom_instruction_master_multi_dataa),
      .A_ci_multi_datab                      (cpu_2_custom_instruction_master_multi_datab),
      .A_ci_multi_done                       (cpu_2_custom_instruction_master_multi_done),
      .A_ci_multi_estatus                    (cpu_2_custom_instruction_master_multi_estatus),
      .A_ci_multi_ipending                   (cpu_2_custom_instruction_master_multi_ipending),
      .A_ci_multi_n                          (cpu_2_custom_instruction_master_multi_n),
      .A_ci_multi_readra                     (cpu_2_custom_instruction_master_multi_readra),
      .A_ci_multi_readrb                     (cpu_2_custom_instruction_master_multi_readrb),
      .A_ci_multi_reset                      (cpu_2_custom_instruction_master_multi_reset),
      .A_ci_multi_result                     (cpu_2_custom_instruction_master_multi_result),
      .A_ci_multi_start                      (cpu_2_custom_instruction_master_multi_start),
      .A_ci_multi_status                     (cpu_2_custom_instruction_master_multi_status),
      .A_ci_multi_writerc                    (cpu_2_custom_instruction_master_multi_writerc),
      .clk                                   (sys_clk),
      .d_address                             (cpu_2_data_master_address),
      .d_byteenable                          (cpu_2_data_master_byteenable),
      .d_irq                                 (cpu_2_data_master_irq),
      .d_read                                (cpu_2_data_master_read),
      .d_readdata                            (cpu_2_data_master_readdata),
      .d_readdatavalid                       (cpu_2_data_master_readdatavalid),
      .d_waitrequest                         (cpu_2_data_master_waitrequest),
      .d_write                               (cpu_2_data_master_write),
      .d_writedata                           (cpu_2_data_master_writedata),
      .i_address                             (cpu_2_instruction_master_address),
      .i_read                                (cpu_2_instruction_master_read),
      .i_readdata                            (cpu_2_instruction_master_readdata),
      .i_readdatavalid                       (cpu_2_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_2_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_2_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_2_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_2_jtag_debug_module_byteenable),
      .jtag_debug_module_debugaccess         (cpu_2_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_2_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_2_jtag_debug_module_readdata),
      .jtag_debug_module_resetrequest        (cpu_2_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_2_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_2_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_2_jtag_debug_module_writedata),
      .reset_n                               (cpu_2_custom_instruction_master_reset_n)
    );

  cpu_2_altera_nios_custom_instr_floating_point_inst_s1_arbitrator the_cpu_2_altera_nios_custom_instr_floating_point_inst_s1
    (
      .clk                                                                                         (sys_clk),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_clk_en                                (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_clk_en),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_dataa                                 (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_dataa),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_datab                                 (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_datab),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done                                  (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa                          (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_n                                     (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_n),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_reset                                 (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_reset),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result                                (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa                        (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select                                (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_select),
      .cpu_2_altera_nios_custom_instr_floating_point_inst_s1_start                                 (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_start),
      .cpu_2_custom_instruction_master_multi_clk_en                                                (cpu_2_custom_instruction_master_multi_clk_en),
      .cpu_2_custom_instruction_master_multi_dataa                                                 (cpu_2_custom_instruction_master_multi_dataa),
      .cpu_2_custom_instruction_master_multi_datab                                                 (cpu_2_custom_instruction_master_multi_datab),
      .cpu_2_custom_instruction_master_multi_n                                                     (cpu_2_custom_instruction_master_multi_n),
      .cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1 (cpu_2_custom_instruction_master_start_cpu_2_altera_nios_custom_instr_floating_point_inst_s1),
      .reset_n                                                                                     (sys_clk_reset_n)
    );

  cpu_2_altera_nios_custom_instr_floating_point_inst the_cpu_2_altera_nios_custom_instr_floating_point_inst
    (
      .clk    (sys_clk),
      .clk_en (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_clk_en),
      .dataa  (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_dataa),
      .datab  (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_datab),
      .done   (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_done),
      .n      (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_n),
      .reset  (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_reset),
      .result (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_result),
      .start  (cpu_2_altera_nios_custom_instr_floating_point_inst_s1_start)
    );

  cpu_3_jtag_debug_module_arbitrator the_cpu_3_jtag_debug_module
    (
      .clk                                                                              (sys_clk),
      .cpu_3_data_master_address_to_slave                                               (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_byteenable                                                     (cpu_3_data_master_byteenable),
      .cpu_3_data_master_debugaccess                                                    (cpu_3_data_master_debugaccess),
      .cpu_3_data_master_granted_cpu_3_jtag_debug_module                                (cpu_3_data_master_granted_cpu_3_jtag_debug_module),
      .cpu_3_data_master_latency_counter                                                (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module                      (cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module),
      .cpu_3_data_master_read                                                           (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module                        (cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_cpu_3_jtag_debug_module                               (cpu_3_data_master_requests_cpu_3_jtag_debug_module),
      .cpu_3_data_master_write                                                          (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                                      (cpu_3_data_master_writedata),
      .cpu_3_instruction_master_address_to_slave                                        (cpu_3_instruction_master_address_to_slave),
      .cpu_3_instruction_master_granted_cpu_3_jtag_debug_module                         (cpu_3_instruction_master_granted_cpu_3_jtag_debug_module),
      .cpu_3_instruction_master_latency_counter                                         (cpu_3_instruction_master_latency_counter),
      .cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module               (cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module),
      .cpu_3_instruction_master_read                                                    (cpu_3_instruction_master_read),
      .cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module                 (cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module),
      .cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_instruction_master_requests_cpu_3_jtag_debug_module                        (cpu_3_instruction_master_requests_cpu_3_jtag_debug_module),
      .cpu_3_jtag_debug_module_address                                                  (cpu_3_jtag_debug_module_address),
      .cpu_3_jtag_debug_module_begintransfer                                            (cpu_3_jtag_debug_module_begintransfer),
      .cpu_3_jtag_debug_module_byteenable                                               (cpu_3_jtag_debug_module_byteenable),
      .cpu_3_jtag_debug_module_chipselect                                               (cpu_3_jtag_debug_module_chipselect),
      .cpu_3_jtag_debug_module_debugaccess                                              (cpu_3_jtag_debug_module_debugaccess),
      .cpu_3_jtag_debug_module_readdata                                                 (cpu_3_jtag_debug_module_readdata),
      .cpu_3_jtag_debug_module_readdata_from_sa                                         (cpu_3_jtag_debug_module_readdata_from_sa),
      .cpu_3_jtag_debug_module_resetrequest                                             (cpu_3_jtag_debug_module_resetrequest),
      .cpu_3_jtag_debug_module_resetrequest_from_sa                                     (cpu_3_jtag_debug_module_resetrequest_from_sa),
      .cpu_3_jtag_debug_module_write                                                    (cpu_3_jtag_debug_module_write),
      .cpu_3_jtag_debug_module_writedata                                                (cpu_3_jtag_debug_module_writedata),
      .d1_cpu_3_jtag_debug_module_end_xfer                                              (d1_cpu_3_jtag_debug_module_end_xfer),
      .reset_n                                                                          (sys_clk_reset_n)
    );

  cpu_3_custom_instruction_master_arbitrator the_cpu_3_custom_instruction_master
    (
      .clk                                                                                         (sys_clk),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa                          (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa                        (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select                                (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select),
      .cpu_3_custom_instruction_master_multi_done                                                  (cpu_3_custom_instruction_master_multi_done),
      .cpu_3_custom_instruction_master_multi_result                                                (cpu_3_custom_instruction_master_multi_result),
      .cpu_3_custom_instruction_master_multi_start                                                 (cpu_3_custom_instruction_master_multi_start),
      .cpu_3_custom_instruction_master_reset_n                                                     (cpu_3_custom_instruction_master_reset_n),
      .cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1 (cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1),
      .reset_n                                                                                     (sys_clk_reset_n)
    );

  cpu_3_data_master_arbitrator the_cpu_3_data_master
    (
      .clk                                                                               (sys_clk),
      .cpu_3_data_master_address                                                         (cpu_3_data_master_address),
      .cpu_3_data_master_address_to_slave                                                (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_byteenable                                                      (cpu_3_data_master_byteenable),
      .cpu_3_data_master_byteenable_nios_system_clock_11_in                              (cpu_3_data_master_byteenable_nios_system_clock_11_in),
      .cpu_3_data_master_byteenable_nios_system_clock_7_in                               (cpu_3_data_master_byteenable_nios_system_clock_7_in),
      .cpu_3_data_master_byteenable_sram_0_avalon_sram_slave                             (cpu_3_data_master_byteenable_sram_0_avalon_sram_slave),
      .cpu_3_data_master_dbs_address                                                     (cpu_3_data_master_dbs_address),
      .cpu_3_data_master_dbs_write_16                                                    (cpu_3_data_master_dbs_write_16),
      .cpu_3_data_master_dbs_write_8                                                     (cpu_3_data_master_dbs_write_8),
      .cpu_3_data_master_granted_cpu_3_jtag_debug_module                                 (cpu_3_data_master_granted_cpu_3_jtag_debug_module),
      .cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave                           (cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave),
      .cpu_3_data_master_granted_keys_s1                                                 (cpu_3_data_master_granted_keys_s1),
      .cpu_3_data_master_granted_mailbox_0_s1                                            (cpu_3_data_master_granted_mailbox_0_s1),
      .cpu_3_data_master_granted_mailbox_1_s1                                            (cpu_3_data_master_granted_mailbox_1_s1),
      .cpu_3_data_master_granted_mailbox_2_s1                                            (cpu_3_data_master_granted_mailbox_2_s1),
      .cpu_3_data_master_granted_mailbox_3_s1                                            (cpu_3_data_master_granted_mailbox_3_s1),
      .cpu_3_data_master_granted_nios_system_clock_11_in                                 (cpu_3_data_master_granted_nios_system_clock_11_in),
      .cpu_3_data_master_granted_nios_system_clock_7_in                                  (cpu_3_data_master_granted_nios_system_clock_7_in),
      .cpu_3_data_master_granted_onchip_memory2_0_s1                                     (cpu_3_data_master_granted_onchip_memory2_0_s1),
      .cpu_3_data_master_granted_onchip_memory2_1_s1                                     (cpu_3_data_master_granted_onchip_memory2_1_s1),
      .cpu_3_data_master_granted_onchip_memory2_2_s1                                     (cpu_3_data_master_granted_onchip_memory2_2_s1),
      .cpu_3_data_master_granted_onchip_memory2_3_s1                                     (cpu_3_data_master_granted_onchip_memory2_3_s1),
      .cpu_3_data_master_granted_performance_counter_0_control_slave                     (cpu_3_data_master_granted_performance_counter_0_control_slave),
      .cpu_3_data_master_granted_sram_0_avalon_sram_slave                                (cpu_3_data_master_granted_sram_0_avalon_sram_slave),
      .cpu_3_data_master_granted_sysid_control_slave                                     (cpu_3_data_master_granted_sysid_control_slave),
      .cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave           (cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_3_data_master_irq                                                             (cpu_3_data_master_irq),
      .cpu_3_data_master_latency_counter                                                 (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module                       (cpu_3_data_master_qualified_request_cpu_3_jtag_debug_module),
      .cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave                 (cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave),
      .cpu_3_data_master_qualified_request_keys_s1                                       (cpu_3_data_master_qualified_request_keys_s1),
      .cpu_3_data_master_qualified_request_mailbox_0_s1                                  (cpu_3_data_master_qualified_request_mailbox_0_s1),
      .cpu_3_data_master_qualified_request_mailbox_1_s1                                  (cpu_3_data_master_qualified_request_mailbox_1_s1),
      .cpu_3_data_master_qualified_request_mailbox_2_s1                                  (cpu_3_data_master_qualified_request_mailbox_2_s1),
      .cpu_3_data_master_qualified_request_mailbox_3_s1                                  (cpu_3_data_master_qualified_request_mailbox_3_s1),
      .cpu_3_data_master_qualified_request_nios_system_clock_11_in                       (cpu_3_data_master_qualified_request_nios_system_clock_11_in),
      .cpu_3_data_master_qualified_request_nios_system_clock_7_in                        (cpu_3_data_master_qualified_request_nios_system_clock_7_in),
      .cpu_3_data_master_qualified_request_onchip_memory2_0_s1                           (cpu_3_data_master_qualified_request_onchip_memory2_0_s1),
      .cpu_3_data_master_qualified_request_onchip_memory2_1_s1                           (cpu_3_data_master_qualified_request_onchip_memory2_1_s1),
      .cpu_3_data_master_qualified_request_onchip_memory2_2_s1                           (cpu_3_data_master_qualified_request_onchip_memory2_2_s1),
      .cpu_3_data_master_qualified_request_onchip_memory2_3_s1                           (cpu_3_data_master_qualified_request_onchip_memory2_3_s1),
      .cpu_3_data_master_qualified_request_performance_counter_0_control_slave           (cpu_3_data_master_qualified_request_performance_counter_0_control_slave),
      .cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave                      (cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_3_data_master_qualified_request_sysid_control_slave                           (cpu_3_data_master_qualified_request_sysid_control_slave),
      .cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave (cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_3_data_master_read                                                            (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module                         (cpu_3_data_master_read_data_valid_cpu_3_jtag_debug_module),
      .cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave                   (cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave),
      .cpu_3_data_master_read_data_valid_keys_s1                                         (cpu_3_data_master_read_data_valid_keys_s1),
      .cpu_3_data_master_read_data_valid_mailbox_0_s1                                    (cpu_3_data_master_read_data_valid_mailbox_0_s1),
      .cpu_3_data_master_read_data_valid_mailbox_1_s1                                    (cpu_3_data_master_read_data_valid_mailbox_1_s1),
      .cpu_3_data_master_read_data_valid_mailbox_2_s1                                    (cpu_3_data_master_read_data_valid_mailbox_2_s1),
      .cpu_3_data_master_read_data_valid_mailbox_3_s1                                    (cpu_3_data_master_read_data_valid_mailbox_3_s1),
      .cpu_3_data_master_read_data_valid_nios_system_clock_11_in                         (cpu_3_data_master_read_data_valid_nios_system_clock_11_in),
      .cpu_3_data_master_read_data_valid_nios_system_clock_7_in                          (cpu_3_data_master_read_data_valid_nios_system_clock_7_in),
      .cpu_3_data_master_read_data_valid_onchip_memory2_0_s1                             (cpu_3_data_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_3_data_master_read_data_valid_onchip_memory2_1_s1                             (cpu_3_data_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_3_data_master_read_data_valid_onchip_memory2_2_s1                             (cpu_3_data_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_3_data_master_read_data_valid_onchip_memory2_3_s1                             (cpu_3_data_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_3_data_master_read_data_valid_performance_counter_0_control_slave             (cpu_3_data_master_read_data_valid_performance_counter_0_control_slave),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave                        (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register         (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_read_data_valid_sysid_control_slave                             (cpu_3_data_master_read_data_valid_sysid_control_slave),
      .cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave   (cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_3_data_master_readdata                                                        (cpu_3_data_master_readdata),
      .cpu_3_data_master_readdatavalid                                                   (cpu_3_data_master_readdatavalid),
      .cpu_3_data_master_requests_cpu_3_jtag_debug_module                                (cpu_3_data_master_requests_cpu_3_jtag_debug_module),
      .cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave                          (cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave),
      .cpu_3_data_master_requests_keys_s1                                                (cpu_3_data_master_requests_keys_s1),
      .cpu_3_data_master_requests_mailbox_0_s1                                           (cpu_3_data_master_requests_mailbox_0_s1),
      .cpu_3_data_master_requests_mailbox_1_s1                                           (cpu_3_data_master_requests_mailbox_1_s1),
      .cpu_3_data_master_requests_mailbox_2_s1                                           (cpu_3_data_master_requests_mailbox_2_s1),
      .cpu_3_data_master_requests_mailbox_3_s1                                           (cpu_3_data_master_requests_mailbox_3_s1),
      .cpu_3_data_master_requests_nios_system_clock_11_in                                (cpu_3_data_master_requests_nios_system_clock_11_in),
      .cpu_3_data_master_requests_nios_system_clock_7_in                                 (cpu_3_data_master_requests_nios_system_clock_7_in),
      .cpu_3_data_master_requests_onchip_memory2_0_s1                                    (cpu_3_data_master_requests_onchip_memory2_0_s1),
      .cpu_3_data_master_requests_onchip_memory2_1_s1                                    (cpu_3_data_master_requests_onchip_memory2_1_s1),
      .cpu_3_data_master_requests_onchip_memory2_2_s1                                    (cpu_3_data_master_requests_onchip_memory2_2_s1),
      .cpu_3_data_master_requests_onchip_memory2_3_s1                                    (cpu_3_data_master_requests_onchip_memory2_3_s1),
      .cpu_3_data_master_requests_performance_counter_0_control_slave                    (cpu_3_data_master_requests_performance_counter_0_control_slave),
      .cpu_3_data_master_requests_sram_0_avalon_sram_slave                               (cpu_3_data_master_requests_sram_0_avalon_sram_slave),
      .cpu_3_data_master_requests_sysid_control_slave                                    (cpu_3_data_master_requests_sysid_control_slave),
      .cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave          (cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_3_data_master_waitrequest                                                     (cpu_3_data_master_waitrequest),
      .cpu_3_data_master_write                                                           (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                                       (cpu_3_data_master_writedata),
      .cpu_3_jtag_debug_module_readdata_from_sa                                          (cpu_3_jtag_debug_module_readdata_from_sa),
      .d1_cpu_3_jtag_debug_module_end_xfer                                               (d1_cpu_3_jtag_debug_module_end_xfer),
      .d1_jtag_uart_3_avalon_jtag_slave_end_xfer                                         (d1_jtag_uart_3_avalon_jtag_slave_end_xfer),
      .d1_keys_s1_end_xfer                                                               (d1_keys_s1_end_xfer),
      .d1_mailbox_0_s1_end_xfer                                                          (d1_mailbox_0_s1_end_xfer),
      .d1_mailbox_1_s1_end_xfer                                                          (d1_mailbox_1_s1_end_xfer),
      .d1_mailbox_2_s1_end_xfer                                                          (d1_mailbox_2_s1_end_xfer),
      .d1_mailbox_3_s1_end_xfer                                                          (d1_mailbox_3_s1_end_xfer),
      .d1_nios_system_clock_11_in_end_xfer                                               (d1_nios_system_clock_11_in_end_xfer),
      .d1_nios_system_clock_7_in_end_xfer                                                (d1_nios_system_clock_7_in_end_xfer),
      .d1_onchip_memory2_0_s1_end_xfer                                                   (d1_onchip_memory2_0_s1_end_xfer),
      .d1_onchip_memory2_1_s1_end_xfer                                                   (d1_onchip_memory2_1_s1_end_xfer),
      .d1_onchip_memory2_2_s1_end_xfer                                                   (d1_onchip_memory2_2_s1_end_xfer),
      .d1_onchip_memory2_3_s1_end_xfer                                                   (d1_onchip_memory2_3_s1_end_xfer),
      .d1_performance_counter_0_control_slave_end_xfer                                   (d1_performance_counter_0_control_slave_end_xfer),
      .d1_sram_0_avalon_sram_slave_end_xfer                                              (d1_sram_0_avalon_sram_slave_end_xfer),
      .d1_sysid_control_slave_end_xfer                                                   (d1_sysid_control_slave_end_xfer),
      .d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer                         (d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer),
      .jtag_uart_3_avalon_jtag_slave_irq_from_sa                                         (jtag_uart_3_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_3_avalon_jtag_slave_readdata_from_sa                                    (jtag_uart_3_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa                                 (jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa),
      .keys_s1_readdata_from_sa                                                          (keys_s1_readdata_from_sa),
      .mailbox_0_s1_readdata_from_sa                                                     (mailbox_0_s1_readdata_from_sa),
      .mailbox_1_s1_readdata_from_sa                                                     (mailbox_1_s1_readdata_from_sa),
      .mailbox_2_s1_readdata_from_sa                                                     (mailbox_2_s1_readdata_from_sa),
      .mailbox_3_s1_readdata_from_sa                                                     (mailbox_3_s1_readdata_from_sa),
      .nios_system_clock_11_in_readdata_from_sa                                          (nios_system_clock_11_in_readdata_from_sa),
      .nios_system_clock_11_in_waitrequest_from_sa                                       (nios_system_clock_11_in_waitrequest_from_sa),
      .nios_system_clock_7_in_readdata_from_sa                                           (nios_system_clock_7_in_readdata_from_sa),
      .nios_system_clock_7_in_waitrequest_from_sa                                        (nios_system_clock_7_in_waitrequest_from_sa),
      .onchip_memory2_0_s1_readdata_from_sa                                              (onchip_memory2_0_s1_readdata_from_sa),
      .onchip_memory2_1_s1_readdata_from_sa                                              (onchip_memory2_1_s1_readdata_from_sa),
      .onchip_memory2_2_s1_readdata_from_sa                                              (onchip_memory2_2_s1_readdata_from_sa),
      .onchip_memory2_3_s1_readdata_from_sa                                              (onchip_memory2_3_s1_readdata_from_sa),
      .performance_counter_0_control_slave_readdata_from_sa                              (performance_counter_0_control_slave_readdata_from_sa),
      .reset_n                                                                           (sys_clk_reset_n),
      .sram_0_avalon_sram_slave_readdata_from_sa                                         (sram_0_avalon_sram_slave_readdata_from_sa),
      .sysid_control_slave_readdata_from_sa                                              (sysid_control_slave_readdata_from_sa),
      .video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa                    (video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa)
    );

  cpu_3_instruction_master_arbitrator the_cpu_3_instruction_master
    (
      .clk                                                                              (sys_clk),
      .cpu_3_instruction_master_address                                                 (cpu_3_instruction_master_address),
      .cpu_3_instruction_master_address_to_slave                                        (cpu_3_instruction_master_address_to_slave),
      .cpu_3_instruction_master_dbs_address                                             (cpu_3_instruction_master_dbs_address),
      .cpu_3_instruction_master_granted_cpu_3_jtag_debug_module                         (cpu_3_instruction_master_granted_cpu_3_jtag_debug_module),
      .cpu_3_instruction_master_granted_nios_system_clock_6_in                          (cpu_3_instruction_master_granted_nios_system_clock_6_in),
      .cpu_3_instruction_master_granted_onchip_memory2_0_s1                             (cpu_3_instruction_master_granted_onchip_memory2_0_s1),
      .cpu_3_instruction_master_granted_onchip_memory2_1_s1                             (cpu_3_instruction_master_granted_onchip_memory2_1_s1),
      .cpu_3_instruction_master_granted_onchip_memory2_2_s1                             (cpu_3_instruction_master_granted_onchip_memory2_2_s1),
      .cpu_3_instruction_master_granted_onchip_memory2_3_s1                             (cpu_3_instruction_master_granted_onchip_memory2_3_s1),
      .cpu_3_instruction_master_granted_sram_0_avalon_sram_slave                        (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave),
      .cpu_3_instruction_master_latency_counter                                         (cpu_3_instruction_master_latency_counter),
      .cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module               (cpu_3_instruction_master_qualified_request_cpu_3_jtag_debug_module),
      .cpu_3_instruction_master_qualified_request_nios_system_clock_6_in                (cpu_3_instruction_master_qualified_request_nios_system_clock_6_in),
      .cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1                   (cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1),
      .cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1                   (cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1),
      .cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1                   (cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1),
      .cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1                   (cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1),
      .cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave              (cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_3_instruction_master_read                                                    (cpu_3_instruction_master_read),
      .cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module                 (cpu_3_instruction_master_read_data_valid_cpu_3_jtag_debug_module),
      .cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in                  (cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in),
      .cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1                     (cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1                     (cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1                     (cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1                     (cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave                (cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_instruction_master_readdata                                                (cpu_3_instruction_master_readdata),
      .cpu_3_instruction_master_readdatavalid                                           (cpu_3_instruction_master_readdatavalid),
      .cpu_3_instruction_master_requests_cpu_3_jtag_debug_module                        (cpu_3_instruction_master_requests_cpu_3_jtag_debug_module),
      .cpu_3_instruction_master_requests_nios_system_clock_6_in                         (cpu_3_instruction_master_requests_nios_system_clock_6_in),
      .cpu_3_instruction_master_requests_onchip_memory2_0_s1                            (cpu_3_instruction_master_requests_onchip_memory2_0_s1),
      .cpu_3_instruction_master_requests_onchip_memory2_1_s1                            (cpu_3_instruction_master_requests_onchip_memory2_1_s1),
      .cpu_3_instruction_master_requests_onchip_memory2_2_s1                            (cpu_3_instruction_master_requests_onchip_memory2_2_s1),
      .cpu_3_instruction_master_requests_onchip_memory2_3_s1                            (cpu_3_instruction_master_requests_onchip_memory2_3_s1),
      .cpu_3_instruction_master_requests_sram_0_avalon_sram_slave                       (cpu_3_instruction_master_requests_sram_0_avalon_sram_slave),
      .cpu_3_instruction_master_waitrequest                                             (cpu_3_instruction_master_waitrequest),
      .cpu_3_jtag_debug_module_readdata_from_sa                                         (cpu_3_jtag_debug_module_readdata_from_sa),
      .d1_cpu_3_jtag_debug_module_end_xfer                                              (d1_cpu_3_jtag_debug_module_end_xfer),
      .d1_nios_system_clock_6_in_end_xfer                                               (d1_nios_system_clock_6_in_end_xfer),
      .d1_onchip_memory2_0_s1_end_xfer                                                  (d1_onchip_memory2_0_s1_end_xfer),
      .d1_onchip_memory2_1_s1_end_xfer                                                  (d1_onchip_memory2_1_s1_end_xfer),
      .d1_onchip_memory2_2_s1_end_xfer                                                  (d1_onchip_memory2_2_s1_end_xfer),
      .d1_onchip_memory2_3_s1_end_xfer                                                  (d1_onchip_memory2_3_s1_end_xfer),
      .d1_sram_0_avalon_sram_slave_end_xfer                                             (d1_sram_0_avalon_sram_slave_end_xfer),
      .nios_system_clock_6_in_readdata_from_sa                                          (nios_system_clock_6_in_readdata_from_sa),
      .nios_system_clock_6_in_waitrequest_from_sa                                       (nios_system_clock_6_in_waitrequest_from_sa),
      .onchip_memory2_0_s1_readdata_from_sa                                             (onchip_memory2_0_s1_readdata_from_sa),
      .onchip_memory2_1_s1_readdata_from_sa                                             (onchip_memory2_1_s1_readdata_from_sa),
      .onchip_memory2_2_s1_readdata_from_sa                                             (onchip_memory2_2_s1_readdata_from_sa),
      .onchip_memory2_3_s1_readdata_from_sa                                             (onchip_memory2_3_s1_readdata_from_sa),
      .reset_n                                                                          (sys_clk_reset_n),
      .sram_0_avalon_sram_slave_readdata_from_sa                                        (sram_0_avalon_sram_slave_readdata_from_sa)
    );

  cpu_3 the_cpu_3
    (
      .A_ci_multi_a                          (cpu_3_custom_instruction_master_multi_a),
      .A_ci_multi_b                          (cpu_3_custom_instruction_master_multi_b),
      .A_ci_multi_c                          (cpu_3_custom_instruction_master_multi_c),
      .A_ci_multi_clk_en                     (cpu_3_custom_instruction_master_multi_clk_en),
      .A_ci_multi_clock                      (cpu_3_custom_instruction_master_multi_clk),
      .A_ci_multi_dataa                      (cpu_3_custom_instruction_master_multi_dataa),
      .A_ci_multi_datab                      (cpu_3_custom_instruction_master_multi_datab),
      .A_ci_multi_done                       (cpu_3_custom_instruction_master_multi_done),
      .A_ci_multi_estatus                    (cpu_3_custom_instruction_master_multi_estatus),
      .A_ci_multi_ipending                   (cpu_3_custom_instruction_master_multi_ipending),
      .A_ci_multi_n                          (cpu_3_custom_instruction_master_multi_n),
      .A_ci_multi_readra                     (cpu_3_custom_instruction_master_multi_readra),
      .A_ci_multi_readrb                     (cpu_3_custom_instruction_master_multi_readrb),
      .A_ci_multi_reset                      (cpu_3_custom_instruction_master_multi_reset),
      .A_ci_multi_result                     (cpu_3_custom_instruction_master_multi_result),
      .A_ci_multi_start                      (cpu_3_custom_instruction_master_multi_start),
      .A_ci_multi_status                     (cpu_3_custom_instruction_master_multi_status),
      .A_ci_multi_writerc                    (cpu_3_custom_instruction_master_multi_writerc),
      .clk                                   (sys_clk),
      .d_address                             (cpu_3_data_master_address),
      .d_byteenable                          (cpu_3_data_master_byteenable),
      .d_irq                                 (cpu_3_data_master_irq),
      .d_read                                (cpu_3_data_master_read),
      .d_readdata                            (cpu_3_data_master_readdata),
      .d_readdatavalid                       (cpu_3_data_master_readdatavalid),
      .d_waitrequest                         (cpu_3_data_master_waitrequest),
      .d_write                               (cpu_3_data_master_write),
      .d_writedata                           (cpu_3_data_master_writedata),
      .i_address                             (cpu_3_instruction_master_address),
      .i_read                                (cpu_3_instruction_master_read),
      .i_readdata                            (cpu_3_instruction_master_readdata),
      .i_readdatavalid                       (cpu_3_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_3_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_3_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_3_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_3_jtag_debug_module_byteenable),
      .jtag_debug_module_debugaccess         (cpu_3_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_3_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_3_jtag_debug_module_readdata),
      .jtag_debug_module_resetrequest        (cpu_3_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_3_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_3_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_3_jtag_debug_module_writedata),
      .reset_n                               (cpu_3_custom_instruction_master_reset_n)
    );

  cpu_3_altera_nios_custom_instr_floating_point_inst_s1_arbitrator the_cpu_3_altera_nios_custom_instr_floating_point_inst_s1
    (
      .clk                                                                                         (sys_clk),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_clk_en                                (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_clk_en),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_dataa                                 (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_dataa),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_datab                                 (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_datab),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done                                  (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa                          (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done_from_sa),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_n                                     (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_n),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_reset                                 (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_reset),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result                                (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa                        (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result_from_sa),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select                                (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_select),
      .cpu_3_altera_nios_custom_instr_floating_point_inst_s1_start                                 (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_start),
      .cpu_3_custom_instruction_master_multi_clk_en                                                (cpu_3_custom_instruction_master_multi_clk_en),
      .cpu_3_custom_instruction_master_multi_dataa                                                 (cpu_3_custom_instruction_master_multi_dataa),
      .cpu_3_custom_instruction_master_multi_datab                                                 (cpu_3_custom_instruction_master_multi_datab),
      .cpu_3_custom_instruction_master_multi_n                                                     (cpu_3_custom_instruction_master_multi_n),
      .cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1 (cpu_3_custom_instruction_master_start_cpu_3_altera_nios_custom_instr_floating_point_inst_s1),
      .reset_n                                                                                     (sys_clk_reset_n)
    );

  cpu_3_altera_nios_custom_instr_floating_point_inst the_cpu_3_altera_nios_custom_instr_floating_point_inst
    (
      .clk    (sys_clk),
      .clk_en (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_clk_en),
      .dataa  (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_dataa),
      .datab  (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_datab),
      .done   (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_done),
      .n      (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_n),
      .reset  (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_reset),
      .result (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_result),
      .start  (cpu_3_altera_nios_custom_instr_floating_point_inst_s1_start)
    );

  jtag_uart_0_avalon_jtag_slave_arbitrator the_jtag_uart_0_avalon_jtag_slave
    (
      .clk                                                                       (sys_clk),
      .cpu_0_data_master_address_to_slave                                        (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave                   (cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_latency_counter                                         (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave         (cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_read                                                    (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave           (cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave                  (cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_write                                                   (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                               (cpu_0_data_master_writedata),
      .d1_jtag_uart_0_avalon_jtag_slave_end_xfer                                 (d1_jtag_uart_0_avalon_jtag_slave_end_xfer),
      .jtag_uart_0_avalon_jtag_slave_address                                     (jtag_uart_0_avalon_jtag_slave_address),
      .jtag_uart_0_avalon_jtag_slave_chipselect                                  (jtag_uart_0_avalon_jtag_slave_chipselect),
      .jtag_uart_0_avalon_jtag_slave_dataavailable                               (jtag_uart_0_avalon_jtag_slave_dataavailable),
      .jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa                       (jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_0_avalon_jtag_slave_irq                                         (jtag_uart_0_avalon_jtag_slave_irq),
      .jtag_uart_0_avalon_jtag_slave_irq_from_sa                                 (jtag_uart_0_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_0_avalon_jtag_slave_read_n                                      (jtag_uart_0_avalon_jtag_slave_read_n),
      .jtag_uart_0_avalon_jtag_slave_readdata                                    (jtag_uart_0_avalon_jtag_slave_readdata),
      .jtag_uart_0_avalon_jtag_slave_readdata_from_sa                            (jtag_uart_0_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_0_avalon_jtag_slave_readyfordata                                (jtag_uart_0_avalon_jtag_slave_readyfordata),
      .jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa                        (jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_0_avalon_jtag_slave_reset_n                                     (jtag_uart_0_avalon_jtag_slave_reset_n),
      .jtag_uart_0_avalon_jtag_slave_waitrequest                                 (jtag_uart_0_avalon_jtag_slave_waitrequest),
      .jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa                         (jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_0_avalon_jtag_slave_write_n                                     (jtag_uart_0_avalon_jtag_slave_write_n),
      .jtag_uart_0_avalon_jtag_slave_writedata                                   (jtag_uart_0_avalon_jtag_slave_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  jtag_uart_0 the_jtag_uart_0
    (
      .av_address     (jtag_uart_0_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_0_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_0_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_0_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_0_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_0_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_0_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_0_avalon_jtag_slave_writedata),
      .clk            (sys_clk),
      .dataavailable  (jtag_uart_0_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_0_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_0_avalon_jtag_slave_reset_n)
    );

  jtag_uart_1_avalon_jtag_slave_arbitrator the_jtag_uart_1_avalon_jtag_slave
    (
      .clk                                                                       (sys_clk),
      .cpu_1_data_master_address_to_slave                                        (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave                   (cpu_1_data_master_granted_jtag_uart_1_avalon_jtag_slave),
      .cpu_1_data_master_latency_counter                                         (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave         (cpu_1_data_master_qualified_request_jtag_uart_1_avalon_jtag_slave),
      .cpu_1_data_master_read                                                    (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave           (cpu_1_data_master_read_data_valid_jtag_uart_1_avalon_jtag_slave),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave                  (cpu_1_data_master_requests_jtag_uart_1_avalon_jtag_slave),
      .cpu_1_data_master_write                                                   (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                               (cpu_1_data_master_writedata),
      .d1_jtag_uart_1_avalon_jtag_slave_end_xfer                                 (d1_jtag_uart_1_avalon_jtag_slave_end_xfer),
      .jtag_uart_1_avalon_jtag_slave_address                                     (jtag_uart_1_avalon_jtag_slave_address),
      .jtag_uart_1_avalon_jtag_slave_chipselect                                  (jtag_uart_1_avalon_jtag_slave_chipselect),
      .jtag_uart_1_avalon_jtag_slave_dataavailable                               (jtag_uart_1_avalon_jtag_slave_dataavailable),
      .jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa                       (jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_1_avalon_jtag_slave_irq                                         (jtag_uart_1_avalon_jtag_slave_irq),
      .jtag_uart_1_avalon_jtag_slave_irq_from_sa                                 (jtag_uart_1_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_1_avalon_jtag_slave_read_n                                      (jtag_uart_1_avalon_jtag_slave_read_n),
      .jtag_uart_1_avalon_jtag_slave_readdata                                    (jtag_uart_1_avalon_jtag_slave_readdata),
      .jtag_uart_1_avalon_jtag_slave_readdata_from_sa                            (jtag_uart_1_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_1_avalon_jtag_slave_readyfordata                                (jtag_uart_1_avalon_jtag_slave_readyfordata),
      .jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa                        (jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_1_avalon_jtag_slave_reset_n                                     (jtag_uart_1_avalon_jtag_slave_reset_n),
      .jtag_uart_1_avalon_jtag_slave_waitrequest                                 (jtag_uart_1_avalon_jtag_slave_waitrequest),
      .jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa                         (jtag_uart_1_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_1_avalon_jtag_slave_write_n                                     (jtag_uart_1_avalon_jtag_slave_write_n),
      .jtag_uart_1_avalon_jtag_slave_writedata                                   (jtag_uart_1_avalon_jtag_slave_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  jtag_uart_1 the_jtag_uart_1
    (
      .av_address     (jtag_uart_1_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_1_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_1_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_1_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_1_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_1_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_1_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_1_avalon_jtag_slave_writedata),
      .clk            (sys_clk),
      .dataavailable  (jtag_uart_1_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_1_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_1_avalon_jtag_slave_reset_n)
    );

  jtag_uart_2_avalon_jtag_slave_arbitrator the_jtag_uart_2_avalon_jtag_slave
    (
      .clk                                                                       (sys_clk),
      .cpu_2_data_master_address_to_slave                                        (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave                   (cpu_2_data_master_granted_jtag_uart_2_avalon_jtag_slave),
      .cpu_2_data_master_latency_counter                                         (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave         (cpu_2_data_master_qualified_request_jtag_uart_2_avalon_jtag_slave),
      .cpu_2_data_master_read                                                    (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave           (cpu_2_data_master_read_data_valid_jtag_uart_2_avalon_jtag_slave),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave                  (cpu_2_data_master_requests_jtag_uart_2_avalon_jtag_slave),
      .cpu_2_data_master_write                                                   (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                               (cpu_2_data_master_writedata),
      .d1_jtag_uart_2_avalon_jtag_slave_end_xfer                                 (d1_jtag_uart_2_avalon_jtag_slave_end_xfer),
      .jtag_uart_2_avalon_jtag_slave_address                                     (jtag_uart_2_avalon_jtag_slave_address),
      .jtag_uart_2_avalon_jtag_slave_chipselect                                  (jtag_uart_2_avalon_jtag_slave_chipselect),
      .jtag_uart_2_avalon_jtag_slave_dataavailable                               (jtag_uart_2_avalon_jtag_slave_dataavailable),
      .jtag_uart_2_avalon_jtag_slave_dataavailable_from_sa                       (jtag_uart_2_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_2_avalon_jtag_slave_irq                                         (jtag_uart_2_avalon_jtag_slave_irq),
      .jtag_uart_2_avalon_jtag_slave_irq_from_sa                                 (jtag_uart_2_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_2_avalon_jtag_slave_read_n                                      (jtag_uart_2_avalon_jtag_slave_read_n),
      .jtag_uart_2_avalon_jtag_slave_readdata                                    (jtag_uart_2_avalon_jtag_slave_readdata),
      .jtag_uart_2_avalon_jtag_slave_readdata_from_sa                            (jtag_uart_2_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_2_avalon_jtag_slave_readyfordata                                (jtag_uart_2_avalon_jtag_slave_readyfordata),
      .jtag_uart_2_avalon_jtag_slave_readyfordata_from_sa                        (jtag_uart_2_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_2_avalon_jtag_slave_reset_n                                     (jtag_uart_2_avalon_jtag_slave_reset_n),
      .jtag_uart_2_avalon_jtag_slave_waitrequest                                 (jtag_uart_2_avalon_jtag_slave_waitrequest),
      .jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa                         (jtag_uart_2_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_2_avalon_jtag_slave_write_n                                     (jtag_uart_2_avalon_jtag_slave_write_n),
      .jtag_uart_2_avalon_jtag_slave_writedata                                   (jtag_uart_2_avalon_jtag_slave_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  jtag_uart_2 the_jtag_uart_2
    (
      .av_address     (jtag_uart_2_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_2_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_2_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_2_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_2_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_2_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_2_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_2_avalon_jtag_slave_writedata),
      .clk            (sys_clk),
      .dataavailable  (jtag_uart_2_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_2_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_2_avalon_jtag_slave_reset_n)
    );

  jtag_uart_3_avalon_jtag_slave_arbitrator the_jtag_uart_3_avalon_jtag_slave
    (
      .clk                                                                       (sys_clk),
      .cpu_3_data_master_address_to_slave                                        (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave                   (cpu_3_data_master_granted_jtag_uart_3_avalon_jtag_slave),
      .cpu_3_data_master_latency_counter                                         (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave         (cpu_3_data_master_qualified_request_jtag_uart_3_avalon_jtag_slave),
      .cpu_3_data_master_read                                                    (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave           (cpu_3_data_master_read_data_valid_jtag_uart_3_avalon_jtag_slave),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave                  (cpu_3_data_master_requests_jtag_uart_3_avalon_jtag_slave),
      .cpu_3_data_master_write                                                   (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                               (cpu_3_data_master_writedata),
      .d1_jtag_uart_3_avalon_jtag_slave_end_xfer                                 (d1_jtag_uart_3_avalon_jtag_slave_end_xfer),
      .jtag_uart_3_avalon_jtag_slave_address                                     (jtag_uart_3_avalon_jtag_slave_address),
      .jtag_uart_3_avalon_jtag_slave_chipselect                                  (jtag_uart_3_avalon_jtag_slave_chipselect),
      .jtag_uart_3_avalon_jtag_slave_dataavailable                               (jtag_uart_3_avalon_jtag_slave_dataavailable),
      .jtag_uart_3_avalon_jtag_slave_dataavailable_from_sa                       (jtag_uart_3_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_3_avalon_jtag_slave_irq                                         (jtag_uart_3_avalon_jtag_slave_irq),
      .jtag_uart_3_avalon_jtag_slave_irq_from_sa                                 (jtag_uart_3_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_3_avalon_jtag_slave_read_n                                      (jtag_uart_3_avalon_jtag_slave_read_n),
      .jtag_uart_3_avalon_jtag_slave_readdata                                    (jtag_uart_3_avalon_jtag_slave_readdata),
      .jtag_uart_3_avalon_jtag_slave_readdata_from_sa                            (jtag_uart_3_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_3_avalon_jtag_slave_readyfordata                                (jtag_uart_3_avalon_jtag_slave_readyfordata),
      .jtag_uart_3_avalon_jtag_slave_readyfordata_from_sa                        (jtag_uart_3_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_3_avalon_jtag_slave_reset_n                                     (jtag_uart_3_avalon_jtag_slave_reset_n),
      .jtag_uart_3_avalon_jtag_slave_waitrequest                                 (jtag_uart_3_avalon_jtag_slave_waitrequest),
      .jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa                         (jtag_uart_3_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_3_avalon_jtag_slave_write_n                                     (jtag_uart_3_avalon_jtag_slave_write_n),
      .jtag_uart_3_avalon_jtag_slave_writedata                                   (jtag_uart_3_avalon_jtag_slave_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  jtag_uart_3 the_jtag_uart_3
    (
      .av_address     (jtag_uart_3_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_3_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_3_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_3_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_3_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_3_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_3_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_3_avalon_jtag_slave_writedata),
      .clk            (sys_clk),
      .dataavailable  (jtag_uart_3_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_3_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_3_avalon_jtag_slave_reset_n)
    );

  keys_s1_arbitrator the_keys_s1
    (
      .clk                                                                       (sys_clk),
      .cpu_0_data_master_address_to_slave                                        (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_keys_s1                                         (cpu_0_data_master_granted_keys_s1),
      .cpu_0_data_master_latency_counter                                         (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_keys_s1                               (cpu_0_data_master_qualified_request_keys_s1),
      .cpu_0_data_master_read                                                    (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_keys_s1                                 (cpu_0_data_master_read_data_valid_keys_s1),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_keys_s1                                        (cpu_0_data_master_requests_keys_s1),
      .cpu_0_data_master_write                                                   (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                               (cpu_0_data_master_writedata),
      .cpu_1_data_master_address_to_slave                                        (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_granted_keys_s1                                         (cpu_1_data_master_granted_keys_s1),
      .cpu_1_data_master_latency_counter                                         (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_keys_s1                               (cpu_1_data_master_qualified_request_keys_s1),
      .cpu_1_data_master_read                                                    (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_keys_s1                                 (cpu_1_data_master_read_data_valid_keys_s1),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_keys_s1                                        (cpu_1_data_master_requests_keys_s1),
      .cpu_1_data_master_write                                                   (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                               (cpu_1_data_master_writedata),
      .cpu_2_data_master_address_to_slave                                        (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_granted_keys_s1                                         (cpu_2_data_master_granted_keys_s1),
      .cpu_2_data_master_latency_counter                                         (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_keys_s1                               (cpu_2_data_master_qualified_request_keys_s1),
      .cpu_2_data_master_read                                                    (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_keys_s1                                 (cpu_2_data_master_read_data_valid_keys_s1),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_keys_s1                                        (cpu_2_data_master_requests_keys_s1),
      .cpu_2_data_master_write                                                   (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                               (cpu_2_data_master_writedata),
      .cpu_3_data_master_address_to_slave                                        (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_granted_keys_s1                                         (cpu_3_data_master_granted_keys_s1),
      .cpu_3_data_master_latency_counter                                         (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_keys_s1                               (cpu_3_data_master_qualified_request_keys_s1),
      .cpu_3_data_master_read                                                    (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_keys_s1                                 (cpu_3_data_master_read_data_valid_keys_s1),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_keys_s1                                        (cpu_3_data_master_requests_keys_s1),
      .cpu_3_data_master_write                                                   (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                               (cpu_3_data_master_writedata),
      .d1_keys_s1_end_xfer                                                       (d1_keys_s1_end_xfer),
      .keys_s1_address                                                           (keys_s1_address),
      .keys_s1_chipselect                                                        (keys_s1_chipselect),
      .keys_s1_readdata                                                          (keys_s1_readdata),
      .keys_s1_readdata_from_sa                                                  (keys_s1_readdata_from_sa),
      .keys_s1_reset_n                                                           (keys_s1_reset_n),
      .keys_s1_write_n                                                           (keys_s1_write_n),
      .keys_s1_writedata                                                         (keys_s1_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  keys the_keys
    (
      .address    (keys_s1_address),
      .chipselect (keys_s1_chipselect),
      .clk        (sys_clk),
      .in_port    (in_port_to_the_keys),
      .readdata   (keys_s1_readdata),
      .reset_n    (keys_s1_reset_n),
      .write_n    (keys_s1_write_n),
      .writedata  (keys_s1_writedata)
    );

  mailbox_0_s1_arbitrator the_mailbox_0_s1
    (
      .clk                                                                       (sys_clk),
      .cpu_0_data_master_address_to_slave                                        (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_mailbox_0_s1                                    (cpu_0_data_master_granted_mailbox_0_s1),
      .cpu_0_data_master_latency_counter                                         (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_mailbox_0_s1                          (cpu_0_data_master_qualified_request_mailbox_0_s1),
      .cpu_0_data_master_read                                                    (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_mailbox_0_s1                            (cpu_0_data_master_read_data_valid_mailbox_0_s1),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_mailbox_0_s1                                   (cpu_0_data_master_requests_mailbox_0_s1),
      .cpu_0_data_master_write                                                   (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                               (cpu_0_data_master_writedata),
      .cpu_1_data_master_address_to_slave                                        (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_granted_mailbox_0_s1                                    (cpu_1_data_master_granted_mailbox_0_s1),
      .cpu_1_data_master_latency_counter                                         (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_mailbox_0_s1                          (cpu_1_data_master_qualified_request_mailbox_0_s1),
      .cpu_1_data_master_read                                                    (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_mailbox_0_s1                            (cpu_1_data_master_read_data_valid_mailbox_0_s1),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_mailbox_0_s1                                   (cpu_1_data_master_requests_mailbox_0_s1),
      .cpu_1_data_master_write                                                   (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                               (cpu_1_data_master_writedata),
      .cpu_2_data_master_address_to_slave                                        (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_granted_mailbox_0_s1                                    (cpu_2_data_master_granted_mailbox_0_s1),
      .cpu_2_data_master_latency_counter                                         (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_mailbox_0_s1                          (cpu_2_data_master_qualified_request_mailbox_0_s1),
      .cpu_2_data_master_read                                                    (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_mailbox_0_s1                            (cpu_2_data_master_read_data_valid_mailbox_0_s1),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_mailbox_0_s1                                   (cpu_2_data_master_requests_mailbox_0_s1),
      .cpu_2_data_master_write                                                   (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                               (cpu_2_data_master_writedata),
      .cpu_3_data_master_address_to_slave                                        (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_granted_mailbox_0_s1                                    (cpu_3_data_master_granted_mailbox_0_s1),
      .cpu_3_data_master_latency_counter                                         (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_mailbox_0_s1                          (cpu_3_data_master_qualified_request_mailbox_0_s1),
      .cpu_3_data_master_read                                                    (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_mailbox_0_s1                            (cpu_3_data_master_read_data_valid_mailbox_0_s1),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_mailbox_0_s1                                   (cpu_3_data_master_requests_mailbox_0_s1),
      .cpu_3_data_master_write                                                   (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                               (cpu_3_data_master_writedata),
      .d1_mailbox_0_s1_end_xfer                                                  (d1_mailbox_0_s1_end_xfer),
      .mailbox_0_s1_address                                                      (mailbox_0_s1_address),
      .mailbox_0_s1_chipselect                                                   (mailbox_0_s1_chipselect),
      .mailbox_0_s1_read                                                         (mailbox_0_s1_read),
      .mailbox_0_s1_readdata                                                     (mailbox_0_s1_readdata),
      .mailbox_0_s1_readdata_from_sa                                             (mailbox_0_s1_readdata_from_sa),
      .mailbox_0_s1_reset_n                                                      (mailbox_0_s1_reset_n),
      .mailbox_0_s1_write                                                        (mailbox_0_s1_write),
      .mailbox_0_s1_writedata                                                    (mailbox_0_s1_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  mailbox_0 the_mailbox_0
    (
      .address       (mailbox_0_s1_address),
      .chipselect    (mailbox_0_s1_chipselect),
      .clk           (sys_clk),
      .data_from_cpu (mailbox_0_s1_writedata),
      .data_to_cpu   (mailbox_0_s1_readdata),
      .read          (mailbox_0_s1_read),
      .reset_n       (mailbox_0_s1_reset_n),
      .write         (mailbox_0_s1_write)
    );

  mailbox_1_s1_arbitrator the_mailbox_1_s1
    (
      .clk                                                                       (sys_clk),
      .cpu_0_data_master_address_to_slave                                        (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_mailbox_1_s1                                    (cpu_0_data_master_granted_mailbox_1_s1),
      .cpu_0_data_master_latency_counter                                         (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_mailbox_1_s1                          (cpu_0_data_master_qualified_request_mailbox_1_s1),
      .cpu_0_data_master_read                                                    (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_mailbox_1_s1                            (cpu_0_data_master_read_data_valid_mailbox_1_s1),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_mailbox_1_s1                                   (cpu_0_data_master_requests_mailbox_1_s1),
      .cpu_0_data_master_write                                                   (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                               (cpu_0_data_master_writedata),
      .cpu_1_data_master_address_to_slave                                        (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_granted_mailbox_1_s1                                    (cpu_1_data_master_granted_mailbox_1_s1),
      .cpu_1_data_master_latency_counter                                         (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_mailbox_1_s1                          (cpu_1_data_master_qualified_request_mailbox_1_s1),
      .cpu_1_data_master_read                                                    (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_mailbox_1_s1                            (cpu_1_data_master_read_data_valid_mailbox_1_s1),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_mailbox_1_s1                                   (cpu_1_data_master_requests_mailbox_1_s1),
      .cpu_1_data_master_write                                                   (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                               (cpu_1_data_master_writedata),
      .cpu_2_data_master_address_to_slave                                        (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_granted_mailbox_1_s1                                    (cpu_2_data_master_granted_mailbox_1_s1),
      .cpu_2_data_master_latency_counter                                         (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_mailbox_1_s1                          (cpu_2_data_master_qualified_request_mailbox_1_s1),
      .cpu_2_data_master_read                                                    (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_mailbox_1_s1                            (cpu_2_data_master_read_data_valid_mailbox_1_s1),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_mailbox_1_s1                                   (cpu_2_data_master_requests_mailbox_1_s1),
      .cpu_2_data_master_write                                                   (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                               (cpu_2_data_master_writedata),
      .cpu_3_data_master_address_to_slave                                        (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_granted_mailbox_1_s1                                    (cpu_3_data_master_granted_mailbox_1_s1),
      .cpu_3_data_master_latency_counter                                         (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_mailbox_1_s1                          (cpu_3_data_master_qualified_request_mailbox_1_s1),
      .cpu_3_data_master_read                                                    (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_mailbox_1_s1                            (cpu_3_data_master_read_data_valid_mailbox_1_s1),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_mailbox_1_s1                                   (cpu_3_data_master_requests_mailbox_1_s1),
      .cpu_3_data_master_write                                                   (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                               (cpu_3_data_master_writedata),
      .d1_mailbox_1_s1_end_xfer                                                  (d1_mailbox_1_s1_end_xfer),
      .mailbox_1_s1_address                                                      (mailbox_1_s1_address),
      .mailbox_1_s1_chipselect                                                   (mailbox_1_s1_chipselect),
      .mailbox_1_s1_read                                                         (mailbox_1_s1_read),
      .mailbox_1_s1_readdata                                                     (mailbox_1_s1_readdata),
      .mailbox_1_s1_readdata_from_sa                                             (mailbox_1_s1_readdata_from_sa),
      .mailbox_1_s1_reset_n                                                      (mailbox_1_s1_reset_n),
      .mailbox_1_s1_write                                                        (mailbox_1_s1_write),
      .mailbox_1_s1_writedata                                                    (mailbox_1_s1_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  mailbox_1 the_mailbox_1
    (
      .address       (mailbox_1_s1_address),
      .chipselect    (mailbox_1_s1_chipselect),
      .clk           (sys_clk),
      .data_from_cpu (mailbox_1_s1_writedata),
      .data_to_cpu   (mailbox_1_s1_readdata),
      .read          (mailbox_1_s1_read),
      .reset_n       (mailbox_1_s1_reset_n),
      .write         (mailbox_1_s1_write)
    );

  mailbox_2_s1_arbitrator the_mailbox_2_s1
    (
      .clk                                                                       (sys_clk),
      .cpu_0_data_master_address_to_slave                                        (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_mailbox_2_s1                                    (cpu_0_data_master_granted_mailbox_2_s1),
      .cpu_0_data_master_latency_counter                                         (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_mailbox_2_s1                          (cpu_0_data_master_qualified_request_mailbox_2_s1),
      .cpu_0_data_master_read                                                    (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_mailbox_2_s1                            (cpu_0_data_master_read_data_valid_mailbox_2_s1),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_mailbox_2_s1                                   (cpu_0_data_master_requests_mailbox_2_s1),
      .cpu_0_data_master_write                                                   (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                               (cpu_0_data_master_writedata),
      .cpu_1_data_master_address_to_slave                                        (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_granted_mailbox_2_s1                                    (cpu_1_data_master_granted_mailbox_2_s1),
      .cpu_1_data_master_latency_counter                                         (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_mailbox_2_s1                          (cpu_1_data_master_qualified_request_mailbox_2_s1),
      .cpu_1_data_master_read                                                    (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_mailbox_2_s1                            (cpu_1_data_master_read_data_valid_mailbox_2_s1),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_mailbox_2_s1                                   (cpu_1_data_master_requests_mailbox_2_s1),
      .cpu_1_data_master_write                                                   (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                               (cpu_1_data_master_writedata),
      .cpu_2_data_master_address_to_slave                                        (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_granted_mailbox_2_s1                                    (cpu_2_data_master_granted_mailbox_2_s1),
      .cpu_2_data_master_latency_counter                                         (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_mailbox_2_s1                          (cpu_2_data_master_qualified_request_mailbox_2_s1),
      .cpu_2_data_master_read                                                    (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_mailbox_2_s1                            (cpu_2_data_master_read_data_valid_mailbox_2_s1),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_mailbox_2_s1                                   (cpu_2_data_master_requests_mailbox_2_s1),
      .cpu_2_data_master_write                                                   (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                               (cpu_2_data_master_writedata),
      .cpu_3_data_master_address_to_slave                                        (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_granted_mailbox_2_s1                                    (cpu_3_data_master_granted_mailbox_2_s1),
      .cpu_3_data_master_latency_counter                                         (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_mailbox_2_s1                          (cpu_3_data_master_qualified_request_mailbox_2_s1),
      .cpu_3_data_master_read                                                    (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_mailbox_2_s1                            (cpu_3_data_master_read_data_valid_mailbox_2_s1),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_mailbox_2_s1                                   (cpu_3_data_master_requests_mailbox_2_s1),
      .cpu_3_data_master_write                                                   (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                               (cpu_3_data_master_writedata),
      .d1_mailbox_2_s1_end_xfer                                                  (d1_mailbox_2_s1_end_xfer),
      .mailbox_2_s1_address                                                      (mailbox_2_s1_address),
      .mailbox_2_s1_chipselect                                                   (mailbox_2_s1_chipselect),
      .mailbox_2_s1_read                                                         (mailbox_2_s1_read),
      .mailbox_2_s1_readdata                                                     (mailbox_2_s1_readdata),
      .mailbox_2_s1_readdata_from_sa                                             (mailbox_2_s1_readdata_from_sa),
      .mailbox_2_s1_reset_n                                                      (mailbox_2_s1_reset_n),
      .mailbox_2_s1_write                                                        (mailbox_2_s1_write),
      .mailbox_2_s1_writedata                                                    (mailbox_2_s1_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  mailbox_2 the_mailbox_2
    (
      .address       (mailbox_2_s1_address),
      .chipselect    (mailbox_2_s1_chipselect),
      .clk           (sys_clk),
      .data_from_cpu (mailbox_2_s1_writedata),
      .data_to_cpu   (mailbox_2_s1_readdata),
      .read          (mailbox_2_s1_read),
      .reset_n       (mailbox_2_s1_reset_n),
      .write         (mailbox_2_s1_write)
    );

  mailbox_3_s1_arbitrator the_mailbox_3_s1
    (
      .clk                                                                       (sys_clk),
      .cpu_0_data_master_address_to_slave                                        (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_mailbox_3_s1                                    (cpu_0_data_master_granted_mailbox_3_s1),
      .cpu_0_data_master_latency_counter                                         (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_mailbox_3_s1                          (cpu_0_data_master_qualified_request_mailbox_3_s1),
      .cpu_0_data_master_read                                                    (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_mailbox_3_s1                            (cpu_0_data_master_read_data_valid_mailbox_3_s1),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_mailbox_3_s1                                   (cpu_0_data_master_requests_mailbox_3_s1),
      .cpu_0_data_master_write                                                   (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                               (cpu_0_data_master_writedata),
      .cpu_1_data_master_address_to_slave                                        (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_granted_mailbox_3_s1                                    (cpu_1_data_master_granted_mailbox_3_s1),
      .cpu_1_data_master_latency_counter                                         (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_mailbox_3_s1                          (cpu_1_data_master_qualified_request_mailbox_3_s1),
      .cpu_1_data_master_read                                                    (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_mailbox_3_s1                            (cpu_1_data_master_read_data_valid_mailbox_3_s1),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_mailbox_3_s1                                   (cpu_1_data_master_requests_mailbox_3_s1),
      .cpu_1_data_master_write                                                   (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                               (cpu_1_data_master_writedata),
      .cpu_2_data_master_address_to_slave                                        (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_granted_mailbox_3_s1                                    (cpu_2_data_master_granted_mailbox_3_s1),
      .cpu_2_data_master_latency_counter                                         (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_mailbox_3_s1                          (cpu_2_data_master_qualified_request_mailbox_3_s1),
      .cpu_2_data_master_read                                                    (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_mailbox_3_s1                            (cpu_2_data_master_read_data_valid_mailbox_3_s1),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_mailbox_3_s1                                   (cpu_2_data_master_requests_mailbox_3_s1),
      .cpu_2_data_master_write                                                   (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                               (cpu_2_data_master_writedata),
      .cpu_3_data_master_address_to_slave                                        (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_granted_mailbox_3_s1                                    (cpu_3_data_master_granted_mailbox_3_s1),
      .cpu_3_data_master_latency_counter                                         (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_mailbox_3_s1                          (cpu_3_data_master_qualified_request_mailbox_3_s1),
      .cpu_3_data_master_read                                                    (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_mailbox_3_s1                            (cpu_3_data_master_read_data_valid_mailbox_3_s1),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_mailbox_3_s1                                   (cpu_3_data_master_requests_mailbox_3_s1),
      .cpu_3_data_master_write                                                   (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                               (cpu_3_data_master_writedata),
      .d1_mailbox_3_s1_end_xfer                                                  (d1_mailbox_3_s1_end_xfer),
      .mailbox_3_s1_address                                                      (mailbox_3_s1_address),
      .mailbox_3_s1_chipselect                                                   (mailbox_3_s1_chipselect),
      .mailbox_3_s1_read                                                         (mailbox_3_s1_read),
      .mailbox_3_s1_readdata                                                     (mailbox_3_s1_readdata),
      .mailbox_3_s1_readdata_from_sa                                             (mailbox_3_s1_readdata_from_sa),
      .mailbox_3_s1_reset_n                                                      (mailbox_3_s1_reset_n),
      .mailbox_3_s1_write                                                        (mailbox_3_s1_write),
      .mailbox_3_s1_writedata                                                    (mailbox_3_s1_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  mailbox_3 the_mailbox_3
    (
      .address       (mailbox_3_s1_address),
      .chipselect    (mailbox_3_s1_chipselect),
      .clk           (sys_clk),
      .data_from_cpu (mailbox_3_s1_writedata),
      .data_to_cpu   (mailbox_3_s1_readdata),
      .read          (mailbox_3_s1_read),
      .reset_n       (mailbox_3_s1_reset_n),
      .write         (mailbox_3_s1_write)
    );

  nios_system_clock_0_in_arbitrator the_nios_system_clock_0_in
    (
      .clk                                                                              (sys_clk),
      .cpu_1_instruction_master_address_to_slave                                        (cpu_1_instruction_master_address_to_slave),
      .cpu_1_instruction_master_dbs_address                                             (cpu_1_instruction_master_dbs_address),
      .cpu_1_instruction_master_granted_nios_system_clock_0_in                          (cpu_1_instruction_master_granted_nios_system_clock_0_in),
      .cpu_1_instruction_master_latency_counter                                         (cpu_1_instruction_master_latency_counter),
      .cpu_1_instruction_master_qualified_request_nios_system_clock_0_in                (cpu_1_instruction_master_qualified_request_nios_system_clock_0_in),
      .cpu_1_instruction_master_read                                                    (cpu_1_instruction_master_read),
      .cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in                  (cpu_1_instruction_master_read_data_valid_nios_system_clock_0_in),
      .cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_instruction_master_requests_nios_system_clock_0_in                         (cpu_1_instruction_master_requests_nios_system_clock_0_in),
      .d1_nios_system_clock_0_in_end_xfer                                               (d1_nios_system_clock_0_in_end_xfer),
      .nios_system_clock_0_in_address                                                   (nios_system_clock_0_in_address),
      .nios_system_clock_0_in_byteenable                                                (nios_system_clock_0_in_byteenable),
      .nios_system_clock_0_in_endofpacket                                               (nios_system_clock_0_in_endofpacket),
      .nios_system_clock_0_in_endofpacket_from_sa                                       (nios_system_clock_0_in_endofpacket_from_sa),
      .nios_system_clock_0_in_nativeaddress                                             (nios_system_clock_0_in_nativeaddress),
      .nios_system_clock_0_in_read                                                      (nios_system_clock_0_in_read),
      .nios_system_clock_0_in_readdata                                                  (nios_system_clock_0_in_readdata),
      .nios_system_clock_0_in_readdata_from_sa                                          (nios_system_clock_0_in_readdata_from_sa),
      .nios_system_clock_0_in_reset_n                                                   (nios_system_clock_0_in_reset_n),
      .nios_system_clock_0_in_waitrequest                                               (nios_system_clock_0_in_waitrequest),
      .nios_system_clock_0_in_waitrequest_from_sa                                       (nios_system_clock_0_in_waitrequest_from_sa),
      .nios_system_clock_0_in_write                                                     (nios_system_clock_0_in_write),
      .reset_n                                                                          (sys_clk_reset_n)
    );

  nios_system_clock_0_out_arbitrator the_nios_system_clock_0_out
    (
      .clk                                                               (sdram_clk),
      .d1_sdram_0_s1_end_xfer                                            (d1_sdram_0_s1_end_xfer),
      .nios_system_clock_0_out_address                                   (nios_system_clock_0_out_address),
      .nios_system_clock_0_out_address_to_slave                          (nios_system_clock_0_out_address_to_slave),
      .nios_system_clock_0_out_byteenable                                (nios_system_clock_0_out_byteenable),
      .nios_system_clock_0_out_granted_sdram_0_s1                        (nios_system_clock_0_out_granted_sdram_0_s1),
      .nios_system_clock_0_out_qualified_request_sdram_0_s1              (nios_system_clock_0_out_qualified_request_sdram_0_s1),
      .nios_system_clock_0_out_read                                      (nios_system_clock_0_out_read),
      .nios_system_clock_0_out_read_data_valid_sdram_0_s1                (nios_system_clock_0_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_0_out_readdata                                  (nios_system_clock_0_out_readdata),
      .nios_system_clock_0_out_requests_sdram_0_s1                       (nios_system_clock_0_out_requests_sdram_0_s1),
      .nios_system_clock_0_out_reset_n                                   (nios_system_clock_0_out_reset_n),
      .nios_system_clock_0_out_waitrequest                               (nios_system_clock_0_out_waitrequest),
      .nios_system_clock_0_out_write                                     (nios_system_clock_0_out_write),
      .nios_system_clock_0_out_writedata                                 (nios_system_clock_0_out_writedata),
      .reset_n                                                           (sdram_clk_reset_n),
      .sdram_0_s1_readdata_from_sa                                       (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_waitrequest_from_sa                                    (sdram_0_s1_waitrequest_from_sa)
    );

  nios_system_clock_0 the_nios_system_clock_0
    (
      .master_address       (nios_system_clock_0_out_address),
      .master_byteenable    (nios_system_clock_0_out_byteenable),
      .master_clk           (sdram_clk),
      .master_endofpacket   (nios_system_clock_0_out_endofpacket),
      .master_nativeaddress (nios_system_clock_0_out_nativeaddress),
      .master_read          (nios_system_clock_0_out_read),
      .master_readdata      (nios_system_clock_0_out_readdata),
      .master_reset_n       (nios_system_clock_0_out_reset_n),
      .master_waitrequest   (nios_system_clock_0_out_waitrequest),
      .master_write         (nios_system_clock_0_out_write),
      .master_writedata     (nios_system_clock_0_out_writedata),
      .slave_address        (nios_system_clock_0_in_address),
      .slave_byteenable     (nios_system_clock_0_in_byteenable),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_0_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_0_in_nativeaddress),
      .slave_read           (nios_system_clock_0_in_read),
      .slave_readdata       (nios_system_clock_0_in_readdata),
      .slave_reset_n        (nios_system_clock_0_in_reset_n),
      .slave_waitrequest    (nios_system_clock_0_in_waitrequest),
      .slave_write          (nios_system_clock_0_in_write),
      .slave_writedata      (nios_system_clock_0_in_writedata)
    );

  nios_system_clock_1_in_arbitrator the_nios_system_clock_1_in
    (
      .clk                                                                       (sys_clk),
      .cpu_1_data_master_address_to_slave                                        (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_byteenable                                              (cpu_1_data_master_byteenable),
      .cpu_1_data_master_byteenable_nios_system_clock_1_in                       (cpu_1_data_master_byteenable_nios_system_clock_1_in),
      .cpu_1_data_master_dbs_address                                             (cpu_1_data_master_dbs_address),
      .cpu_1_data_master_dbs_write_16                                            (cpu_1_data_master_dbs_write_16),
      .cpu_1_data_master_granted_nios_system_clock_1_in                          (cpu_1_data_master_granted_nios_system_clock_1_in),
      .cpu_1_data_master_latency_counter                                         (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_nios_system_clock_1_in                (cpu_1_data_master_qualified_request_nios_system_clock_1_in),
      .cpu_1_data_master_read                                                    (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_nios_system_clock_1_in                  (cpu_1_data_master_read_data_valid_nios_system_clock_1_in),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_nios_system_clock_1_in                         (cpu_1_data_master_requests_nios_system_clock_1_in),
      .cpu_1_data_master_write                                                   (cpu_1_data_master_write),
      .d1_nios_system_clock_1_in_end_xfer                                        (d1_nios_system_clock_1_in_end_xfer),
      .nios_system_clock_1_in_address                                            (nios_system_clock_1_in_address),
      .nios_system_clock_1_in_byteenable                                         (nios_system_clock_1_in_byteenable),
      .nios_system_clock_1_in_endofpacket                                        (nios_system_clock_1_in_endofpacket),
      .nios_system_clock_1_in_endofpacket_from_sa                                (nios_system_clock_1_in_endofpacket_from_sa),
      .nios_system_clock_1_in_nativeaddress                                      (nios_system_clock_1_in_nativeaddress),
      .nios_system_clock_1_in_read                                               (nios_system_clock_1_in_read),
      .nios_system_clock_1_in_readdata                                           (nios_system_clock_1_in_readdata),
      .nios_system_clock_1_in_readdata_from_sa                                   (nios_system_clock_1_in_readdata_from_sa),
      .nios_system_clock_1_in_reset_n                                            (nios_system_clock_1_in_reset_n),
      .nios_system_clock_1_in_waitrequest                                        (nios_system_clock_1_in_waitrequest),
      .nios_system_clock_1_in_waitrequest_from_sa                                (nios_system_clock_1_in_waitrequest_from_sa),
      .nios_system_clock_1_in_write                                              (nios_system_clock_1_in_write),
      .nios_system_clock_1_in_writedata                                          (nios_system_clock_1_in_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  nios_system_clock_1_out_arbitrator the_nios_system_clock_1_out
    (
      .clk                                                               (sdram_clk),
      .d1_sdram_0_s1_end_xfer                                            (d1_sdram_0_s1_end_xfer),
      .nios_system_clock_1_out_address                                   (nios_system_clock_1_out_address),
      .nios_system_clock_1_out_address_to_slave                          (nios_system_clock_1_out_address_to_slave),
      .nios_system_clock_1_out_byteenable                                (nios_system_clock_1_out_byteenable),
      .nios_system_clock_1_out_granted_sdram_0_s1                        (nios_system_clock_1_out_granted_sdram_0_s1),
      .nios_system_clock_1_out_qualified_request_sdram_0_s1              (nios_system_clock_1_out_qualified_request_sdram_0_s1),
      .nios_system_clock_1_out_read                                      (nios_system_clock_1_out_read),
      .nios_system_clock_1_out_read_data_valid_sdram_0_s1                (nios_system_clock_1_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_1_out_readdata                                  (nios_system_clock_1_out_readdata),
      .nios_system_clock_1_out_requests_sdram_0_s1                       (nios_system_clock_1_out_requests_sdram_0_s1),
      .nios_system_clock_1_out_reset_n                                   (nios_system_clock_1_out_reset_n),
      .nios_system_clock_1_out_waitrequest                               (nios_system_clock_1_out_waitrequest),
      .nios_system_clock_1_out_write                                     (nios_system_clock_1_out_write),
      .nios_system_clock_1_out_writedata                                 (nios_system_clock_1_out_writedata),
      .reset_n                                                           (sdram_clk_reset_n),
      .sdram_0_s1_readdata_from_sa                                       (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_waitrequest_from_sa                                    (sdram_0_s1_waitrequest_from_sa)
    );

  nios_system_clock_1 the_nios_system_clock_1
    (
      .master_address       (nios_system_clock_1_out_address),
      .master_byteenable    (nios_system_clock_1_out_byteenable),
      .master_clk           (sdram_clk),
      .master_endofpacket   (nios_system_clock_1_out_endofpacket),
      .master_nativeaddress (nios_system_clock_1_out_nativeaddress),
      .master_read          (nios_system_clock_1_out_read),
      .master_readdata      (nios_system_clock_1_out_readdata),
      .master_reset_n       (nios_system_clock_1_out_reset_n),
      .master_waitrequest   (nios_system_clock_1_out_waitrequest),
      .master_write         (nios_system_clock_1_out_write),
      .master_writedata     (nios_system_clock_1_out_writedata),
      .slave_address        (nios_system_clock_1_in_address),
      .slave_byteenable     (nios_system_clock_1_in_byteenable),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_1_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_1_in_nativeaddress),
      .slave_read           (nios_system_clock_1_in_read),
      .slave_readdata       (nios_system_clock_1_in_readdata),
      .slave_reset_n        (nios_system_clock_1_in_reset_n),
      .slave_waitrequest    (nios_system_clock_1_in_waitrequest),
      .slave_write          (nios_system_clock_1_in_write),
      .slave_writedata      (nios_system_clock_1_in_writedata)
    );

  nios_system_clock_10_in_arbitrator the_nios_system_clock_10_in
    (
      .clk                                                                       (sys_clk),
      .cpu_2_data_master_address_to_slave                                        (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_byteenable                                              (cpu_2_data_master_byteenable),
      .cpu_2_data_master_byteenable_nios_system_clock_10_in                      (cpu_2_data_master_byteenable_nios_system_clock_10_in),
      .cpu_2_data_master_dbs_address                                             (cpu_2_data_master_dbs_address),
      .cpu_2_data_master_dbs_write_8                                             (cpu_2_data_master_dbs_write_8),
      .cpu_2_data_master_granted_nios_system_clock_10_in                         (cpu_2_data_master_granted_nios_system_clock_10_in),
      .cpu_2_data_master_latency_counter                                         (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_nios_system_clock_10_in               (cpu_2_data_master_qualified_request_nios_system_clock_10_in),
      .cpu_2_data_master_read                                                    (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_nios_system_clock_10_in                 (cpu_2_data_master_read_data_valid_nios_system_clock_10_in),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_nios_system_clock_10_in                        (cpu_2_data_master_requests_nios_system_clock_10_in),
      .cpu_2_data_master_write                                                   (cpu_2_data_master_write),
      .d1_nios_system_clock_10_in_end_xfer                                       (d1_nios_system_clock_10_in_end_xfer),
      .nios_system_clock_10_in_address                                           (nios_system_clock_10_in_address),
      .nios_system_clock_10_in_endofpacket                                       (nios_system_clock_10_in_endofpacket),
      .nios_system_clock_10_in_endofpacket_from_sa                               (nios_system_clock_10_in_endofpacket_from_sa),
      .nios_system_clock_10_in_nativeaddress                                     (nios_system_clock_10_in_nativeaddress),
      .nios_system_clock_10_in_read                                              (nios_system_clock_10_in_read),
      .nios_system_clock_10_in_readdata                                          (nios_system_clock_10_in_readdata),
      .nios_system_clock_10_in_readdata_from_sa                                  (nios_system_clock_10_in_readdata_from_sa),
      .nios_system_clock_10_in_reset_n                                           (nios_system_clock_10_in_reset_n),
      .nios_system_clock_10_in_waitrequest                                       (nios_system_clock_10_in_waitrequest),
      .nios_system_clock_10_in_waitrequest_from_sa                               (nios_system_clock_10_in_waitrequest_from_sa),
      .nios_system_clock_10_in_write                                             (nios_system_clock_10_in_write),
      .nios_system_clock_10_in_writedata                                         (nios_system_clock_10_in_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  nios_system_clock_10_out_arbitrator the_nios_system_clock_10_out
    (
      .clk                                                                     (clk_0),
      .clocks_0_avalon_clocks_slave_readdata_from_sa                           (clocks_0_avalon_clocks_slave_readdata_from_sa),
      .d1_clocks_0_avalon_clocks_slave_end_xfer                                (d1_clocks_0_avalon_clocks_slave_end_xfer),
      .nios_system_clock_10_out_address                                        (nios_system_clock_10_out_address),
      .nios_system_clock_10_out_address_to_slave                               (nios_system_clock_10_out_address_to_slave),
      .nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave           (nios_system_clock_10_out_granted_clocks_0_avalon_clocks_slave),
      .nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave (nios_system_clock_10_out_qualified_request_clocks_0_avalon_clocks_slave),
      .nios_system_clock_10_out_read                                           (nios_system_clock_10_out_read),
      .nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave   (nios_system_clock_10_out_read_data_valid_clocks_0_avalon_clocks_slave),
      .nios_system_clock_10_out_readdata                                       (nios_system_clock_10_out_readdata),
      .nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave          (nios_system_clock_10_out_requests_clocks_0_avalon_clocks_slave),
      .nios_system_clock_10_out_reset_n                                        (nios_system_clock_10_out_reset_n),
      .nios_system_clock_10_out_waitrequest                                    (nios_system_clock_10_out_waitrequest),
      .nios_system_clock_10_out_write                                          (nios_system_clock_10_out_write),
      .nios_system_clock_10_out_writedata                                      (nios_system_clock_10_out_writedata),
      .reset_n                                                                 (clk_0_reset_n)
    );

  nios_system_clock_10 the_nios_system_clock_10
    (
      .master_address       (nios_system_clock_10_out_address),
      .master_clk           (clk_0),
      .master_endofpacket   (nios_system_clock_10_out_endofpacket),
      .master_nativeaddress (nios_system_clock_10_out_nativeaddress),
      .master_read          (nios_system_clock_10_out_read),
      .master_readdata      (nios_system_clock_10_out_readdata),
      .master_reset_n       (nios_system_clock_10_out_reset_n),
      .master_waitrequest   (nios_system_clock_10_out_waitrequest),
      .master_write         (nios_system_clock_10_out_write),
      .master_writedata     (nios_system_clock_10_out_writedata),
      .slave_address        (nios_system_clock_10_in_address),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_10_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_10_in_nativeaddress),
      .slave_read           (nios_system_clock_10_in_read),
      .slave_readdata       (nios_system_clock_10_in_readdata),
      .slave_reset_n        (nios_system_clock_10_in_reset_n),
      .slave_waitrequest    (nios_system_clock_10_in_waitrequest),
      .slave_write          (nios_system_clock_10_in_write),
      .slave_writedata      (nios_system_clock_10_in_writedata)
    );

  nios_system_clock_11_in_arbitrator the_nios_system_clock_11_in
    (
      .clk                                                                       (sys_clk),
      .cpu_3_data_master_address_to_slave                                        (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_byteenable                                              (cpu_3_data_master_byteenable),
      .cpu_3_data_master_byteenable_nios_system_clock_11_in                      (cpu_3_data_master_byteenable_nios_system_clock_11_in),
      .cpu_3_data_master_dbs_address                                             (cpu_3_data_master_dbs_address),
      .cpu_3_data_master_dbs_write_8                                             (cpu_3_data_master_dbs_write_8),
      .cpu_3_data_master_granted_nios_system_clock_11_in                         (cpu_3_data_master_granted_nios_system_clock_11_in),
      .cpu_3_data_master_latency_counter                                         (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_nios_system_clock_11_in               (cpu_3_data_master_qualified_request_nios_system_clock_11_in),
      .cpu_3_data_master_read                                                    (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_nios_system_clock_11_in                 (cpu_3_data_master_read_data_valid_nios_system_clock_11_in),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_nios_system_clock_11_in                        (cpu_3_data_master_requests_nios_system_clock_11_in),
      .cpu_3_data_master_write                                                   (cpu_3_data_master_write),
      .d1_nios_system_clock_11_in_end_xfer                                       (d1_nios_system_clock_11_in_end_xfer),
      .nios_system_clock_11_in_address                                           (nios_system_clock_11_in_address),
      .nios_system_clock_11_in_endofpacket                                       (nios_system_clock_11_in_endofpacket),
      .nios_system_clock_11_in_endofpacket_from_sa                               (nios_system_clock_11_in_endofpacket_from_sa),
      .nios_system_clock_11_in_nativeaddress                                     (nios_system_clock_11_in_nativeaddress),
      .nios_system_clock_11_in_read                                              (nios_system_clock_11_in_read),
      .nios_system_clock_11_in_readdata                                          (nios_system_clock_11_in_readdata),
      .nios_system_clock_11_in_readdata_from_sa                                  (nios_system_clock_11_in_readdata_from_sa),
      .nios_system_clock_11_in_reset_n                                           (nios_system_clock_11_in_reset_n),
      .nios_system_clock_11_in_waitrequest                                       (nios_system_clock_11_in_waitrequest),
      .nios_system_clock_11_in_waitrequest_from_sa                               (nios_system_clock_11_in_waitrequest_from_sa),
      .nios_system_clock_11_in_write                                             (nios_system_clock_11_in_write),
      .nios_system_clock_11_in_writedata                                         (nios_system_clock_11_in_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  nios_system_clock_11_out_arbitrator the_nios_system_clock_11_out
    (
      .clk                                                                     (clk_0),
      .clocks_0_avalon_clocks_slave_readdata_from_sa                           (clocks_0_avalon_clocks_slave_readdata_from_sa),
      .d1_clocks_0_avalon_clocks_slave_end_xfer                                (d1_clocks_0_avalon_clocks_slave_end_xfer),
      .nios_system_clock_11_out_address                                        (nios_system_clock_11_out_address),
      .nios_system_clock_11_out_address_to_slave                               (nios_system_clock_11_out_address_to_slave),
      .nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave           (nios_system_clock_11_out_granted_clocks_0_avalon_clocks_slave),
      .nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave (nios_system_clock_11_out_qualified_request_clocks_0_avalon_clocks_slave),
      .nios_system_clock_11_out_read                                           (nios_system_clock_11_out_read),
      .nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave   (nios_system_clock_11_out_read_data_valid_clocks_0_avalon_clocks_slave),
      .nios_system_clock_11_out_readdata                                       (nios_system_clock_11_out_readdata),
      .nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave          (nios_system_clock_11_out_requests_clocks_0_avalon_clocks_slave),
      .nios_system_clock_11_out_reset_n                                        (nios_system_clock_11_out_reset_n),
      .nios_system_clock_11_out_waitrequest                                    (nios_system_clock_11_out_waitrequest),
      .nios_system_clock_11_out_write                                          (nios_system_clock_11_out_write),
      .nios_system_clock_11_out_writedata                                      (nios_system_clock_11_out_writedata),
      .reset_n                                                                 (clk_0_reset_n)
    );

  nios_system_clock_11 the_nios_system_clock_11
    (
      .master_address       (nios_system_clock_11_out_address),
      .master_clk           (clk_0),
      .master_endofpacket   (nios_system_clock_11_out_endofpacket),
      .master_nativeaddress (nios_system_clock_11_out_nativeaddress),
      .master_read          (nios_system_clock_11_out_read),
      .master_readdata      (nios_system_clock_11_out_readdata),
      .master_reset_n       (nios_system_clock_11_out_reset_n),
      .master_waitrequest   (nios_system_clock_11_out_waitrequest),
      .master_write         (nios_system_clock_11_out_write),
      .master_writedata     (nios_system_clock_11_out_writedata),
      .slave_address        (nios_system_clock_11_in_address),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_11_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_11_in_nativeaddress),
      .slave_read           (nios_system_clock_11_in_read),
      .slave_readdata       (nios_system_clock_11_in_readdata),
      .slave_reset_n        (nios_system_clock_11_in_reset_n),
      .slave_waitrequest    (nios_system_clock_11_in_waitrequest),
      .slave_write          (nios_system_clock_11_in_write),
      .slave_writedata      (nios_system_clock_11_in_writedata)
    );

  nios_system_clock_2_in_arbitrator the_nios_system_clock_2_in
    (
      .clk                                                               (sys_clk),
      .cpu_0_instruction_master_address_to_slave                         (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_dbs_address                              (cpu_0_instruction_master_dbs_address),
      .cpu_0_instruction_master_granted_nios_system_clock_2_in           (cpu_0_instruction_master_granted_nios_system_clock_2_in),
      .cpu_0_instruction_master_latency_counter                          (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_nios_system_clock_2_in (cpu_0_instruction_master_qualified_request_nios_system_clock_2_in),
      .cpu_0_instruction_master_read                                     (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in   (cpu_0_instruction_master_read_data_valid_nios_system_clock_2_in),
      .cpu_0_instruction_master_requests_nios_system_clock_2_in          (cpu_0_instruction_master_requests_nios_system_clock_2_in),
      .d1_nios_system_clock_2_in_end_xfer                                (d1_nios_system_clock_2_in_end_xfer),
      .nios_system_clock_2_in_address                                    (nios_system_clock_2_in_address),
      .nios_system_clock_2_in_byteenable                                 (nios_system_clock_2_in_byteenable),
      .nios_system_clock_2_in_endofpacket                                (nios_system_clock_2_in_endofpacket),
      .nios_system_clock_2_in_endofpacket_from_sa                        (nios_system_clock_2_in_endofpacket_from_sa),
      .nios_system_clock_2_in_nativeaddress                              (nios_system_clock_2_in_nativeaddress),
      .nios_system_clock_2_in_read                                       (nios_system_clock_2_in_read),
      .nios_system_clock_2_in_readdata                                   (nios_system_clock_2_in_readdata),
      .nios_system_clock_2_in_readdata_from_sa                           (nios_system_clock_2_in_readdata_from_sa),
      .nios_system_clock_2_in_reset_n                                    (nios_system_clock_2_in_reset_n),
      .nios_system_clock_2_in_waitrequest                                (nios_system_clock_2_in_waitrequest),
      .nios_system_clock_2_in_waitrequest_from_sa                        (nios_system_clock_2_in_waitrequest_from_sa),
      .nios_system_clock_2_in_write                                      (nios_system_clock_2_in_write),
      .reset_n                                                           (sys_clk_reset_n)
    );

  nios_system_clock_2_out_arbitrator the_nios_system_clock_2_out
    (
      .clk                                                               (sdram_clk),
      .d1_sdram_0_s1_end_xfer                                            (d1_sdram_0_s1_end_xfer),
      .nios_system_clock_2_out_address                                   (nios_system_clock_2_out_address),
      .nios_system_clock_2_out_address_to_slave                          (nios_system_clock_2_out_address_to_slave),
      .nios_system_clock_2_out_byteenable                                (nios_system_clock_2_out_byteenable),
      .nios_system_clock_2_out_granted_sdram_0_s1                        (nios_system_clock_2_out_granted_sdram_0_s1),
      .nios_system_clock_2_out_qualified_request_sdram_0_s1              (nios_system_clock_2_out_qualified_request_sdram_0_s1),
      .nios_system_clock_2_out_read                                      (nios_system_clock_2_out_read),
      .nios_system_clock_2_out_read_data_valid_sdram_0_s1                (nios_system_clock_2_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_2_out_readdata                                  (nios_system_clock_2_out_readdata),
      .nios_system_clock_2_out_requests_sdram_0_s1                       (nios_system_clock_2_out_requests_sdram_0_s1),
      .nios_system_clock_2_out_reset_n                                   (nios_system_clock_2_out_reset_n),
      .nios_system_clock_2_out_waitrequest                               (nios_system_clock_2_out_waitrequest),
      .nios_system_clock_2_out_write                                     (nios_system_clock_2_out_write),
      .nios_system_clock_2_out_writedata                                 (nios_system_clock_2_out_writedata),
      .reset_n                                                           (sdram_clk_reset_n),
      .sdram_0_s1_readdata_from_sa                                       (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_waitrequest_from_sa                                    (sdram_0_s1_waitrequest_from_sa)
    );

  nios_system_clock_2 the_nios_system_clock_2
    (
      .master_address       (nios_system_clock_2_out_address),
      .master_byteenable    (nios_system_clock_2_out_byteenable),
      .master_clk           (sdram_clk),
      .master_endofpacket   (nios_system_clock_2_out_endofpacket),
      .master_nativeaddress (nios_system_clock_2_out_nativeaddress),
      .master_read          (nios_system_clock_2_out_read),
      .master_readdata      (nios_system_clock_2_out_readdata),
      .master_reset_n       (nios_system_clock_2_out_reset_n),
      .master_waitrequest   (nios_system_clock_2_out_waitrequest),
      .master_write         (nios_system_clock_2_out_write),
      .master_writedata     (nios_system_clock_2_out_writedata),
      .slave_address        (nios_system_clock_2_in_address),
      .slave_byteenable     (nios_system_clock_2_in_byteenable),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_2_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_2_in_nativeaddress),
      .slave_read           (nios_system_clock_2_in_read),
      .slave_readdata       (nios_system_clock_2_in_readdata),
      .slave_reset_n        (nios_system_clock_2_in_reset_n),
      .slave_waitrequest    (nios_system_clock_2_in_waitrequest),
      .slave_write          (nios_system_clock_2_in_write),
      .slave_writedata      (nios_system_clock_2_in_writedata)
    );

  nios_system_clock_3_in_arbitrator the_nios_system_clock_3_in
    (
      .clk                                                                       (sys_clk),
      .cpu_0_data_master_address_to_slave                                        (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                              (cpu_0_data_master_byteenable),
      .cpu_0_data_master_byteenable_nios_system_clock_3_in                       (cpu_0_data_master_byteenable_nios_system_clock_3_in),
      .cpu_0_data_master_dbs_address                                             (cpu_0_data_master_dbs_address),
      .cpu_0_data_master_dbs_write_16                                            (cpu_0_data_master_dbs_write_16),
      .cpu_0_data_master_granted_nios_system_clock_3_in                          (cpu_0_data_master_granted_nios_system_clock_3_in),
      .cpu_0_data_master_latency_counter                                         (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_nios_system_clock_3_in                (cpu_0_data_master_qualified_request_nios_system_clock_3_in),
      .cpu_0_data_master_read                                                    (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_nios_system_clock_3_in                  (cpu_0_data_master_read_data_valid_nios_system_clock_3_in),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_nios_system_clock_3_in                         (cpu_0_data_master_requests_nios_system_clock_3_in),
      .cpu_0_data_master_write                                                   (cpu_0_data_master_write),
      .d1_nios_system_clock_3_in_end_xfer                                        (d1_nios_system_clock_3_in_end_xfer),
      .nios_system_clock_3_in_address                                            (nios_system_clock_3_in_address),
      .nios_system_clock_3_in_byteenable                                         (nios_system_clock_3_in_byteenable),
      .nios_system_clock_3_in_endofpacket                                        (nios_system_clock_3_in_endofpacket),
      .nios_system_clock_3_in_endofpacket_from_sa                                (nios_system_clock_3_in_endofpacket_from_sa),
      .nios_system_clock_3_in_nativeaddress                                      (nios_system_clock_3_in_nativeaddress),
      .nios_system_clock_3_in_read                                               (nios_system_clock_3_in_read),
      .nios_system_clock_3_in_readdata                                           (nios_system_clock_3_in_readdata),
      .nios_system_clock_3_in_readdata_from_sa                                   (nios_system_clock_3_in_readdata_from_sa),
      .nios_system_clock_3_in_reset_n                                            (nios_system_clock_3_in_reset_n),
      .nios_system_clock_3_in_waitrequest                                        (nios_system_clock_3_in_waitrequest),
      .nios_system_clock_3_in_waitrequest_from_sa                                (nios_system_clock_3_in_waitrequest_from_sa),
      .nios_system_clock_3_in_write                                              (nios_system_clock_3_in_write),
      .nios_system_clock_3_in_writedata                                          (nios_system_clock_3_in_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  nios_system_clock_3_out_arbitrator the_nios_system_clock_3_out
    (
      .clk                                                               (sdram_clk),
      .d1_sdram_0_s1_end_xfer                                            (d1_sdram_0_s1_end_xfer),
      .nios_system_clock_3_out_address                                   (nios_system_clock_3_out_address),
      .nios_system_clock_3_out_address_to_slave                          (nios_system_clock_3_out_address_to_slave),
      .nios_system_clock_3_out_byteenable                                (nios_system_clock_3_out_byteenable),
      .nios_system_clock_3_out_granted_sdram_0_s1                        (nios_system_clock_3_out_granted_sdram_0_s1),
      .nios_system_clock_3_out_qualified_request_sdram_0_s1              (nios_system_clock_3_out_qualified_request_sdram_0_s1),
      .nios_system_clock_3_out_read                                      (nios_system_clock_3_out_read),
      .nios_system_clock_3_out_read_data_valid_sdram_0_s1                (nios_system_clock_3_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_3_out_readdata                                  (nios_system_clock_3_out_readdata),
      .nios_system_clock_3_out_requests_sdram_0_s1                       (nios_system_clock_3_out_requests_sdram_0_s1),
      .nios_system_clock_3_out_reset_n                                   (nios_system_clock_3_out_reset_n),
      .nios_system_clock_3_out_waitrequest                               (nios_system_clock_3_out_waitrequest),
      .nios_system_clock_3_out_write                                     (nios_system_clock_3_out_write),
      .nios_system_clock_3_out_writedata                                 (nios_system_clock_3_out_writedata),
      .reset_n                                                           (sdram_clk_reset_n),
      .sdram_0_s1_readdata_from_sa                                       (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_waitrequest_from_sa                                    (sdram_0_s1_waitrequest_from_sa)
    );

  nios_system_clock_3 the_nios_system_clock_3
    (
      .master_address       (nios_system_clock_3_out_address),
      .master_byteenable    (nios_system_clock_3_out_byteenable),
      .master_clk           (sdram_clk),
      .master_endofpacket   (nios_system_clock_3_out_endofpacket),
      .master_nativeaddress (nios_system_clock_3_out_nativeaddress),
      .master_read          (nios_system_clock_3_out_read),
      .master_readdata      (nios_system_clock_3_out_readdata),
      .master_reset_n       (nios_system_clock_3_out_reset_n),
      .master_waitrequest   (nios_system_clock_3_out_waitrequest),
      .master_write         (nios_system_clock_3_out_write),
      .master_writedata     (nios_system_clock_3_out_writedata),
      .slave_address        (nios_system_clock_3_in_address),
      .slave_byteenable     (nios_system_clock_3_in_byteenable),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_3_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_3_in_nativeaddress),
      .slave_read           (nios_system_clock_3_in_read),
      .slave_readdata       (nios_system_clock_3_in_readdata),
      .slave_reset_n        (nios_system_clock_3_in_reset_n),
      .slave_waitrequest    (nios_system_clock_3_in_waitrequest),
      .slave_write          (nios_system_clock_3_in_write),
      .slave_writedata      (nios_system_clock_3_in_writedata)
    );

  nios_system_clock_4_in_arbitrator the_nios_system_clock_4_in
    (
      .clk                                                                              (sys_clk),
      .cpu_2_instruction_master_address_to_slave                                        (cpu_2_instruction_master_address_to_slave),
      .cpu_2_instruction_master_dbs_address                                             (cpu_2_instruction_master_dbs_address),
      .cpu_2_instruction_master_granted_nios_system_clock_4_in                          (cpu_2_instruction_master_granted_nios_system_clock_4_in),
      .cpu_2_instruction_master_latency_counter                                         (cpu_2_instruction_master_latency_counter),
      .cpu_2_instruction_master_qualified_request_nios_system_clock_4_in                (cpu_2_instruction_master_qualified_request_nios_system_clock_4_in),
      .cpu_2_instruction_master_read                                                    (cpu_2_instruction_master_read),
      .cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in                  (cpu_2_instruction_master_read_data_valid_nios_system_clock_4_in),
      .cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_instruction_master_requests_nios_system_clock_4_in                         (cpu_2_instruction_master_requests_nios_system_clock_4_in),
      .d1_nios_system_clock_4_in_end_xfer                                               (d1_nios_system_clock_4_in_end_xfer),
      .nios_system_clock_4_in_address                                                   (nios_system_clock_4_in_address),
      .nios_system_clock_4_in_byteenable                                                (nios_system_clock_4_in_byteenable),
      .nios_system_clock_4_in_endofpacket                                               (nios_system_clock_4_in_endofpacket),
      .nios_system_clock_4_in_endofpacket_from_sa                                       (nios_system_clock_4_in_endofpacket_from_sa),
      .nios_system_clock_4_in_nativeaddress                                             (nios_system_clock_4_in_nativeaddress),
      .nios_system_clock_4_in_read                                                      (nios_system_clock_4_in_read),
      .nios_system_clock_4_in_readdata                                                  (nios_system_clock_4_in_readdata),
      .nios_system_clock_4_in_readdata_from_sa                                          (nios_system_clock_4_in_readdata_from_sa),
      .nios_system_clock_4_in_reset_n                                                   (nios_system_clock_4_in_reset_n),
      .nios_system_clock_4_in_waitrequest                                               (nios_system_clock_4_in_waitrequest),
      .nios_system_clock_4_in_waitrequest_from_sa                                       (nios_system_clock_4_in_waitrequest_from_sa),
      .nios_system_clock_4_in_write                                                     (nios_system_clock_4_in_write),
      .reset_n                                                                          (sys_clk_reset_n)
    );

  nios_system_clock_4_out_arbitrator the_nios_system_clock_4_out
    (
      .clk                                                               (sdram_clk),
      .d1_sdram_0_s1_end_xfer                                            (d1_sdram_0_s1_end_xfer),
      .nios_system_clock_4_out_address                                   (nios_system_clock_4_out_address),
      .nios_system_clock_4_out_address_to_slave                          (nios_system_clock_4_out_address_to_slave),
      .nios_system_clock_4_out_byteenable                                (nios_system_clock_4_out_byteenable),
      .nios_system_clock_4_out_granted_sdram_0_s1                        (nios_system_clock_4_out_granted_sdram_0_s1),
      .nios_system_clock_4_out_qualified_request_sdram_0_s1              (nios_system_clock_4_out_qualified_request_sdram_0_s1),
      .nios_system_clock_4_out_read                                      (nios_system_clock_4_out_read),
      .nios_system_clock_4_out_read_data_valid_sdram_0_s1                (nios_system_clock_4_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_4_out_readdata                                  (nios_system_clock_4_out_readdata),
      .nios_system_clock_4_out_requests_sdram_0_s1                       (nios_system_clock_4_out_requests_sdram_0_s1),
      .nios_system_clock_4_out_reset_n                                   (nios_system_clock_4_out_reset_n),
      .nios_system_clock_4_out_waitrequest                               (nios_system_clock_4_out_waitrequest),
      .nios_system_clock_4_out_write                                     (nios_system_clock_4_out_write),
      .nios_system_clock_4_out_writedata                                 (nios_system_clock_4_out_writedata),
      .reset_n                                                           (sdram_clk_reset_n),
      .sdram_0_s1_readdata_from_sa                                       (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_waitrequest_from_sa                                    (sdram_0_s1_waitrequest_from_sa)
    );

  nios_system_clock_4 the_nios_system_clock_4
    (
      .master_address       (nios_system_clock_4_out_address),
      .master_byteenable    (nios_system_clock_4_out_byteenable),
      .master_clk           (sdram_clk),
      .master_endofpacket   (nios_system_clock_4_out_endofpacket),
      .master_nativeaddress (nios_system_clock_4_out_nativeaddress),
      .master_read          (nios_system_clock_4_out_read),
      .master_readdata      (nios_system_clock_4_out_readdata),
      .master_reset_n       (nios_system_clock_4_out_reset_n),
      .master_waitrequest   (nios_system_clock_4_out_waitrequest),
      .master_write         (nios_system_clock_4_out_write),
      .master_writedata     (nios_system_clock_4_out_writedata),
      .slave_address        (nios_system_clock_4_in_address),
      .slave_byteenable     (nios_system_clock_4_in_byteenable),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_4_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_4_in_nativeaddress),
      .slave_read           (nios_system_clock_4_in_read),
      .slave_readdata       (nios_system_clock_4_in_readdata),
      .slave_reset_n        (nios_system_clock_4_in_reset_n),
      .slave_waitrequest    (nios_system_clock_4_in_waitrequest),
      .slave_write          (nios_system_clock_4_in_write),
      .slave_writedata      (nios_system_clock_4_in_writedata)
    );

  nios_system_clock_5_in_arbitrator the_nios_system_clock_5_in
    (
      .clk                                                                       (sys_clk),
      .cpu_2_data_master_address_to_slave                                        (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_byteenable                                              (cpu_2_data_master_byteenable),
      .cpu_2_data_master_byteenable_nios_system_clock_5_in                       (cpu_2_data_master_byteenable_nios_system_clock_5_in),
      .cpu_2_data_master_dbs_address                                             (cpu_2_data_master_dbs_address),
      .cpu_2_data_master_dbs_write_16                                            (cpu_2_data_master_dbs_write_16),
      .cpu_2_data_master_granted_nios_system_clock_5_in                          (cpu_2_data_master_granted_nios_system_clock_5_in),
      .cpu_2_data_master_latency_counter                                         (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_nios_system_clock_5_in                (cpu_2_data_master_qualified_request_nios_system_clock_5_in),
      .cpu_2_data_master_read                                                    (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_nios_system_clock_5_in                  (cpu_2_data_master_read_data_valid_nios_system_clock_5_in),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_nios_system_clock_5_in                         (cpu_2_data_master_requests_nios_system_clock_5_in),
      .cpu_2_data_master_write                                                   (cpu_2_data_master_write),
      .d1_nios_system_clock_5_in_end_xfer                                        (d1_nios_system_clock_5_in_end_xfer),
      .nios_system_clock_5_in_address                                            (nios_system_clock_5_in_address),
      .nios_system_clock_5_in_byteenable                                         (nios_system_clock_5_in_byteenable),
      .nios_system_clock_5_in_endofpacket                                        (nios_system_clock_5_in_endofpacket),
      .nios_system_clock_5_in_endofpacket_from_sa                                (nios_system_clock_5_in_endofpacket_from_sa),
      .nios_system_clock_5_in_nativeaddress                                      (nios_system_clock_5_in_nativeaddress),
      .nios_system_clock_5_in_read                                               (nios_system_clock_5_in_read),
      .nios_system_clock_5_in_readdata                                           (nios_system_clock_5_in_readdata),
      .nios_system_clock_5_in_readdata_from_sa                                   (nios_system_clock_5_in_readdata_from_sa),
      .nios_system_clock_5_in_reset_n                                            (nios_system_clock_5_in_reset_n),
      .nios_system_clock_5_in_waitrequest                                        (nios_system_clock_5_in_waitrequest),
      .nios_system_clock_5_in_waitrequest_from_sa                                (nios_system_clock_5_in_waitrequest_from_sa),
      .nios_system_clock_5_in_write                                              (nios_system_clock_5_in_write),
      .nios_system_clock_5_in_writedata                                          (nios_system_clock_5_in_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  nios_system_clock_5_out_arbitrator the_nios_system_clock_5_out
    (
      .clk                                                               (sdram_clk),
      .d1_sdram_0_s1_end_xfer                                            (d1_sdram_0_s1_end_xfer),
      .nios_system_clock_5_out_address                                   (nios_system_clock_5_out_address),
      .nios_system_clock_5_out_address_to_slave                          (nios_system_clock_5_out_address_to_slave),
      .nios_system_clock_5_out_byteenable                                (nios_system_clock_5_out_byteenable),
      .nios_system_clock_5_out_granted_sdram_0_s1                        (nios_system_clock_5_out_granted_sdram_0_s1),
      .nios_system_clock_5_out_qualified_request_sdram_0_s1              (nios_system_clock_5_out_qualified_request_sdram_0_s1),
      .nios_system_clock_5_out_read                                      (nios_system_clock_5_out_read),
      .nios_system_clock_5_out_read_data_valid_sdram_0_s1                (nios_system_clock_5_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_5_out_readdata                                  (nios_system_clock_5_out_readdata),
      .nios_system_clock_5_out_requests_sdram_0_s1                       (nios_system_clock_5_out_requests_sdram_0_s1),
      .nios_system_clock_5_out_reset_n                                   (nios_system_clock_5_out_reset_n),
      .nios_system_clock_5_out_waitrequest                               (nios_system_clock_5_out_waitrequest),
      .nios_system_clock_5_out_write                                     (nios_system_clock_5_out_write),
      .nios_system_clock_5_out_writedata                                 (nios_system_clock_5_out_writedata),
      .reset_n                                                           (sdram_clk_reset_n),
      .sdram_0_s1_readdata_from_sa                                       (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_waitrequest_from_sa                                    (sdram_0_s1_waitrequest_from_sa)
    );

  nios_system_clock_5 the_nios_system_clock_5
    (
      .master_address       (nios_system_clock_5_out_address),
      .master_byteenable    (nios_system_clock_5_out_byteenable),
      .master_clk           (sdram_clk),
      .master_endofpacket   (nios_system_clock_5_out_endofpacket),
      .master_nativeaddress (nios_system_clock_5_out_nativeaddress),
      .master_read          (nios_system_clock_5_out_read),
      .master_readdata      (nios_system_clock_5_out_readdata),
      .master_reset_n       (nios_system_clock_5_out_reset_n),
      .master_waitrequest   (nios_system_clock_5_out_waitrequest),
      .master_write         (nios_system_clock_5_out_write),
      .master_writedata     (nios_system_clock_5_out_writedata),
      .slave_address        (nios_system_clock_5_in_address),
      .slave_byteenable     (nios_system_clock_5_in_byteenable),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_5_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_5_in_nativeaddress),
      .slave_read           (nios_system_clock_5_in_read),
      .slave_readdata       (nios_system_clock_5_in_readdata),
      .slave_reset_n        (nios_system_clock_5_in_reset_n),
      .slave_waitrequest    (nios_system_clock_5_in_waitrequest),
      .slave_write          (nios_system_clock_5_in_write),
      .slave_writedata      (nios_system_clock_5_in_writedata)
    );

  nios_system_clock_6_in_arbitrator the_nios_system_clock_6_in
    (
      .clk                                                                              (sys_clk),
      .cpu_3_instruction_master_address_to_slave                                        (cpu_3_instruction_master_address_to_slave),
      .cpu_3_instruction_master_dbs_address                                             (cpu_3_instruction_master_dbs_address),
      .cpu_3_instruction_master_granted_nios_system_clock_6_in                          (cpu_3_instruction_master_granted_nios_system_clock_6_in),
      .cpu_3_instruction_master_latency_counter                                         (cpu_3_instruction_master_latency_counter),
      .cpu_3_instruction_master_qualified_request_nios_system_clock_6_in                (cpu_3_instruction_master_qualified_request_nios_system_clock_6_in),
      .cpu_3_instruction_master_read                                                    (cpu_3_instruction_master_read),
      .cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in                  (cpu_3_instruction_master_read_data_valid_nios_system_clock_6_in),
      .cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_instruction_master_requests_nios_system_clock_6_in                         (cpu_3_instruction_master_requests_nios_system_clock_6_in),
      .d1_nios_system_clock_6_in_end_xfer                                               (d1_nios_system_clock_6_in_end_xfer),
      .nios_system_clock_6_in_address                                                   (nios_system_clock_6_in_address),
      .nios_system_clock_6_in_byteenable                                                (nios_system_clock_6_in_byteenable),
      .nios_system_clock_6_in_endofpacket                                               (nios_system_clock_6_in_endofpacket),
      .nios_system_clock_6_in_endofpacket_from_sa                                       (nios_system_clock_6_in_endofpacket_from_sa),
      .nios_system_clock_6_in_nativeaddress                                             (nios_system_clock_6_in_nativeaddress),
      .nios_system_clock_6_in_read                                                      (nios_system_clock_6_in_read),
      .nios_system_clock_6_in_readdata                                                  (nios_system_clock_6_in_readdata),
      .nios_system_clock_6_in_readdata_from_sa                                          (nios_system_clock_6_in_readdata_from_sa),
      .nios_system_clock_6_in_reset_n                                                   (nios_system_clock_6_in_reset_n),
      .nios_system_clock_6_in_waitrequest                                               (nios_system_clock_6_in_waitrequest),
      .nios_system_clock_6_in_waitrequest_from_sa                                       (nios_system_clock_6_in_waitrequest_from_sa),
      .nios_system_clock_6_in_write                                                     (nios_system_clock_6_in_write),
      .reset_n                                                                          (sys_clk_reset_n)
    );

  nios_system_clock_6_out_arbitrator the_nios_system_clock_6_out
    (
      .clk                                                               (sdram_clk),
      .d1_sdram_0_s1_end_xfer                                            (d1_sdram_0_s1_end_xfer),
      .nios_system_clock_6_out_address                                   (nios_system_clock_6_out_address),
      .nios_system_clock_6_out_address_to_slave                          (nios_system_clock_6_out_address_to_slave),
      .nios_system_clock_6_out_byteenable                                (nios_system_clock_6_out_byteenable),
      .nios_system_clock_6_out_granted_sdram_0_s1                        (nios_system_clock_6_out_granted_sdram_0_s1),
      .nios_system_clock_6_out_qualified_request_sdram_0_s1              (nios_system_clock_6_out_qualified_request_sdram_0_s1),
      .nios_system_clock_6_out_read                                      (nios_system_clock_6_out_read),
      .nios_system_clock_6_out_read_data_valid_sdram_0_s1                (nios_system_clock_6_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_6_out_readdata                                  (nios_system_clock_6_out_readdata),
      .nios_system_clock_6_out_requests_sdram_0_s1                       (nios_system_clock_6_out_requests_sdram_0_s1),
      .nios_system_clock_6_out_reset_n                                   (nios_system_clock_6_out_reset_n),
      .nios_system_clock_6_out_waitrequest                               (nios_system_clock_6_out_waitrequest),
      .nios_system_clock_6_out_write                                     (nios_system_clock_6_out_write),
      .nios_system_clock_6_out_writedata                                 (nios_system_clock_6_out_writedata),
      .reset_n                                                           (sdram_clk_reset_n),
      .sdram_0_s1_readdata_from_sa                                       (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_waitrequest_from_sa                                    (sdram_0_s1_waitrequest_from_sa)
    );

  nios_system_clock_6 the_nios_system_clock_6
    (
      .master_address       (nios_system_clock_6_out_address),
      .master_byteenable    (nios_system_clock_6_out_byteenable),
      .master_clk           (sdram_clk),
      .master_endofpacket   (nios_system_clock_6_out_endofpacket),
      .master_nativeaddress (nios_system_clock_6_out_nativeaddress),
      .master_read          (nios_system_clock_6_out_read),
      .master_readdata      (nios_system_clock_6_out_readdata),
      .master_reset_n       (nios_system_clock_6_out_reset_n),
      .master_waitrequest   (nios_system_clock_6_out_waitrequest),
      .master_write         (nios_system_clock_6_out_write),
      .master_writedata     (nios_system_clock_6_out_writedata),
      .slave_address        (nios_system_clock_6_in_address),
      .slave_byteenable     (nios_system_clock_6_in_byteenable),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_6_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_6_in_nativeaddress),
      .slave_read           (nios_system_clock_6_in_read),
      .slave_readdata       (nios_system_clock_6_in_readdata),
      .slave_reset_n        (nios_system_clock_6_in_reset_n),
      .slave_waitrequest    (nios_system_clock_6_in_waitrequest),
      .slave_write          (nios_system_clock_6_in_write),
      .slave_writedata      (nios_system_clock_6_in_writedata)
    );

  nios_system_clock_7_in_arbitrator the_nios_system_clock_7_in
    (
      .clk                                                                       (sys_clk),
      .cpu_3_data_master_address_to_slave                                        (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_byteenable                                              (cpu_3_data_master_byteenable),
      .cpu_3_data_master_byteenable_nios_system_clock_7_in                       (cpu_3_data_master_byteenable_nios_system_clock_7_in),
      .cpu_3_data_master_dbs_address                                             (cpu_3_data_master_dbs_address),
      .cpu_3_data_master_dbs_write_16                                            (cpu_3_data_master_dbs_write_16),
      .cpu_3_data_master_granted_nios_system_clock_7_in                          (cpu_3_data_master_granted_nios_system_clock_7_in),
      .cpu_3_data_master_latency_counter                                         (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_nios_system_clock_7_in                (cpu_3_data_master_qualified_request_nios_system_clock_7_in),
      .cpu_3_data_master_read                                                    (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_nios_system_clock_7_in                  (cpu_3_data_master_read_data_valid_nios_system_clock_7_in),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_nios_system_clock_7_in                         (cpu_3_data_master_requests_nios_system_clock_7_in),
      .cpu_3_data_master_write                                                   (cpu_3_data_master_write),
      .d1_nios_system_clock_7_in_end_xfer                                        (d1_nios_system_clock_7_in_end_xfer),
      .nios_system_clock_7_in_address                                            (nios_system_clock_7_in_address),
      .nios_system_clock_7_in_byteenable                                         (nios_system_clock_7_in_byteenable),
      .nios_system_clock_7_in_endofpacket                                        (nios_system_clock_7_in_endofpacket),
      .nios_system_clock_7_in_endofpacket_from_sa                                (nios_system_clock_7_in_endofpacket_from_sa),
      .nios_system_clock_7_in_nativeaddress                                      (nios_system_clock_7_in_nativeaddress),
      .nios_system_clock_7_in_read                                               (nios_system_clock_7_in_read),
      .nios_system_clock_7_in_readdata                                           (nios_system_clock_7_in_readdata),
      .nios_system_clock_7_in_readdata_from_sa                                   (nios_system_clock_7_in_readdata_from_sa),
      .nios_system_clock_7_in_reset_n                                            (nios_system_clock_7_in_reset_n),
      .nios_system_clock_7_in_waitrequest                                        (nios_system_clock_7_in_waitrequest),
      .nios_system_clock_7_in_waitrequest_from_sa                                (nios_system_clock_7_in_waitrequest_from_sa),
      .nios_system_clock_7_in_write                                              (nios_system_clock_7_in_write),
      .nios_system_clock_7_in_writedata                                          (nios_system_clock_7_in_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  nios_system_clock_7_out_arbitrator the_nios_system_clock_7_out
    (
      .clk                                                               (sdram_clk),
      .d1_sdram_0_s1_end_xfer                                            (d1_sdram_0_s1_end_xfer),
      .nios_system_clock_7_out_address                                   (nios_system_clock_7_out_address),
      .nios_system_clock_7_out_address_to_slave                          (nios_system_clock_7_out_address_to_slave),
      .nios_system_clock_7_out_byteenable                                (nios_system_clock_7_out_byteenable),
      .nios_system_clock_7_out_granted_sdram_0_s1                        (nios_system_clock_7_out_granted_sdram_0_s1),
      .nios_system_clock_7_out_qualified_request_sdram_0_s1              (nios_system_clock_7_out_qualified_request_sdram_0_s1),
      .nios_system_clock_7_out_read                                      (nios_system_clock_7_out_read),
      .nios_system_clock_7_out_read_data_valid_sdram_0_s1                (nios_system_clock_7_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_7_out_readdata                                  (nios_system_clock_7_out_readdata),
      .nios_system_clock_7_out_requests_sdram_0_s1                       (nios_system_clock_7_out_requests_sdram_0_s1),
      .nios_system_clock_7_out_reset_n                                   (nios_system_clock_7_out_reset_n),
      .nios_system_clock_7_out_waitrequest                               (nios_system_clock_7_out_waitrequest),
      .nios_system_clock_7_out_write                                     (nios_system_clock_7_out_write),
      .nios_system_clock_7_out_writedata                                 (nios_system_clock_7_out_writedata),
      .reset_n                                                           (sdram_clk_reset_n),
      .sdram_0_s1_readdata_from_sa                                       (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_waitrequest_from_sa                                    (sdram_0_s1_waitrequest_from_sa)
    );

  nios_system_clock_7 the_nios_system_clock_7
    (
      .master_address       (nios_system_clock_7_out_address),
      .master_byteenable    (nios_system_clock_7_out_byteenable),
      .master_clk           (sdram_clk),
      .master_endofpacket   (nios_system_clock_7_out_endofpacket),
      .master_nativeaddress (nios_system_clock_7_out_nativeaddress),
      .master_read          (nios_system_clock_7_out_read),
      .master_readdata      (nios_system_clock_7_out_readdata),
      .master_reset_n       (nios_system_clock_7_out_reset_n),
      .master_waitrequest   (nios_system_clock_7_out_waitrequest),
      .master_write         (nios_system_clock_7_out_write),
      .master_writedata     (nios_system_clock_7_out_writedata),
      .slave_address        (nios_system_clock_7_in_address),
      .slave_byteenable     (nios_system_clock_7_in_byteenable),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_7_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_7_in_nativeaddress),
      .slave_read           (nios_system_clock_7_in_read),
      .slave_readdata       (nios_system_clock_7_in_readdata),
      .slave_reset_n        (nios_system_clock_7_in_reset_n),
      .slave_waitrequest    (nios_system_clock_7_in_waitrequest),
      .slave_write          (nios_system_clock_7_in_write),
      .slave_writedata      (nios_system_clock_7_in_writedata)
    );

  nios_system_clock_8_in_arbitrator the_nios_system_clock_8_in
    (
      .clk                                                                       (sys_clk),
      .cpu_1_data_master_address_to_slave                                        (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_byteenable                                              (cpu_1_data_master_byteenable),
      .cpu_1_data_master_byteenable_nios_system_clock_8_in                       (cpu_1_data_master_byteenable_nios_system_clock_8_in),
      .cpu_1_data_master_dbs_address                                             (cpu_1_data_master_dbs_address),
      .cpu_1_data_master_dbs_write_8                                             (cpu_1_data_master_dbs_write_8),
      .cpu_1_data_master_granted_nios_system_clock_8_in                          (cpu_1_data_master_granted_nios_system_clock_8_in),
      .cpu_1_data_master_latency_counter                                         (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_nios_system_clock_8_in                (cpu_1_data_master_qualified_request_nios_system_clock_8_in),
      .cpu_1_data_master_read                                                    (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_nios_system_clock_8_in                  (cpu_1_data_master_read_data_valid_nios_system_clock_8_in),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_nios_system_clock_8_in                         (cpu_1_data_master_requests_nios_system_clock_8_in),
      .cpu_1_data_master_write                                                   (cpu_1_data_master_write),
      .d1_nios_system_clock_8_in_end_xfer                                        (d1_nios_system_clock_8_in_end_xfer),
      .nios_system_clock_8_in_address                                            (nios_system_clock_8_in_address),
      .nios_system_clock_8_in_endofpacket                                        (nios_system_clock_8_in_endofpacket),
      .nios_system_clock_8_in_endofpacket_from_sa                                (nios_system_clock_8_in_endofpacket_from_sa),
      .nios_system_clock_8_in_nativeaddress                                      (nios_system_clock_8_in_nativeaddress),
      .nios_system_clock_8_in_read                                               (nios_system_clock_8_in_read),
      .nios_system_clock_8_in_readdata                                           (nios_system_clock_8_in_readdata),
      .nios_system_clock_8_in_readdata_from_sa                                   (nios_system_clock_8_in_readdata_from_sa),
      .nios_system_clock_8_in_reset_n                                            (nios_system_clock_8_in_reset_n),
      .nios_system_clock_8_in_waitrequest                                        (nios_system_clock_8_in_waitrequest),
      .nios_system_clock_8_in_waitrequest_from_sa                                (nios_system_clock_8_in_waitrequest_from_sa),
      .nios_system_clock_8_in_write                                              (nios_system_clock_8_in_write),
      .nios_system_clock_8_in_writedata                                          (nios_system_clock_8_in_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  nios_system_clock_8_out_arbitrator the_nios_system_clock_8_out
    (
      .clk                                                                    (clk_0),
      .clocks_0_avalon_clocks_slave_readdata_from_sa                          (clocks_0_avalon_clocks_slave_readdata_from_sa),
      .d1_clocks_0_avalon_clocks_slave_end_xfer                               (d1_clocks_0_avalon_clocks_slave_end_xfer),
      .nios_system_clock_8_out_address                                        (nios_system_clock_8_out_address),
      .nios_system_clock_8_out_address_to_slave                               (nios_system_clock_8_out_address_to_slave),
      .nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave           (nios_system_clock_8_out_granted_clocks_0_avalon_clocks_slave),
      .nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave (nios_system_clock_8_out_qualified_request_clocks_0_avalon_clocks_slave),
      .nios_system_clock_8_out_read                                           (nios_system_clock_8_out_read),
      .nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave   (nios_system_clock_8_out_read_data_valid_clocks_0_avalon_clocks_slave),
      .nios_system_clock_8_out_readdata                                       (nios_system_clock_8_out_readdata),
      .nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave          (nios_system_clock_8_out_requests_clocks_0_avalon_clocks_slave),
      .nios_system_clock_8_out_reset_n                                        (nios_system_clock_8_out_reset_n),
      .nios_system_clock_8_out_waitrequest                                    (nios_system_clock_8_out_waitrequest),
      .nios_system_clock_8_out_write                                          (nios_system_clock_8_out_write),
      .nios_system_clock_8_out_writedata                                      (nios_system_clock_8_out_writedata),
      .reset_n                                                                (clk_0_reset_n)
    );

  nios_system_clock_8 the_nios_system_clock_8
    (
      .master_address       (nios_system_clock_8_out_address),
      .master_clk           (clk_0),
      .master_endofpacket   (nios_system_clock_8_out_endofpacket),
      .master_nativeaddress (nios_system_clock_8_out_nativeaddress),
      .master_read          (nios_system_clock_8_out_read),
      .master_readdata      (nios_system_clock_8_out_readdata),
      .master_reset_n       (nios_system_clock_8_out_reset_n),
      .master_waitrequest   (nios_system_clock_8_out_waitrequest),
      .master_write         (nios_system_clock_8_out_write),
      .master_writedata     (nios_system_clock_8_out_writedata),
      .slave_address        (nios_system_clock_8_in_address),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_8_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_8_in_nativeaddress),
      .slave_read           (nios_system_clock_8_in_read),
      .slave_readdata       (nios_system_clock_8_in_readdata),
      .slave_reset_n        (nios_system_clock_8_in_reset_n),
      .slave_waitrequest    (nios_system_clock_8_in_waitrequest),
      .slave_write          (nios_system_clock_8_in_write),
      .slave_writedata      (nios_system_clock_8_in_writedata)
    );

  nios_system_clock_9_in_arbitrator the_nios_system_clock_9_in
    (
      .clk                                                                       (sys_clk),
      .cpu_0_data_master_address_to_slave                                        (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                              (cpu_0_data_master_byteenable),
      .cpu_0_data_master_byteenable_nios_system_clock_9_in                       (cpu_0_data_master_byteenable_nios_system_clock_9_in),
      .cpu_0_data_master_dbs_address                                             (cpu_0_data_master_dbs_address),
      .cpu_0_data_master_dbs_write_8                                             (cpu_0_data_master_dbs_write_8),
      .cpu_0_data_master_granted_nios_system_clock_9_in                          (cpu_0_data_master_granted_nios_system_clock_9_in),
      .cpu_0_data_master_latency_counter                                         (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_nios_system_clock_9_in                (cpu_0_data_master_qualified_request_nios_system_clock_9_in),
      .cpu_0_data_master_read                                                    (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_nios_system_clock_9_in                  (cpu_0_data_master_read_data_valid_nios_system_clock_9_in),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_nios_system_clock_9_in                         (cpu_0_data_master_requests_nios_system_clock_9_in),
      .cpu_0_data_master_write                                                   (cpu_0_data_master_write),
      .d1_nios_system_clock_9_in_end_xfer                                        (d1_nios_system_clock_9_in_end_xfer),
      .nios_system_clock_9_in_address                                            (nios_system_clock_9_in_address),
      .nios_system_clock_9_in_endofpacket                                        (nios_system_clock_9_in_endofpacket),
      .nios_system_clock_9_in_endofpacket_from_sa                                (nios_system_clock_9_in_endofpacket_from_sa),
      .nios_system_clock_9_in_nativeaddress                                      (nios_system_clock_9_in_nativeaddress),
      .nios_system_clock_9_in_read                                               (nios_system_clock_9_in_read),
      .nios_system_clock_9_in_readdata                                           (nios_system_clock_9_in_readdata),
      .nios_system_clock_9_in_readdata_from_sa                                   (nios_system_clock_9_in_readdata_from_sa),
      .nios_system_clock_9_in_reset_n                                            (nios_system_clock_9_in_reset_n),
      .nios_system_clock_9_in_waitrequest                                        (nios_system_clock_9_in_waitrequest),
      .nios_system_clock_9_in_waitrequest_from_sa                                (nios_system_clock_9_in_waitrequest_from_sa),
      .nios_system_clock_9_in_write                                              (nios_system_clock_9_in_write),
      .nios_system_clock_9_in_writedata                                          (nios_system_clock_9_in_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  nios_system_clock_9_out_arbitrator the_nios_system_clock_9_out
    (
      .clk                                                                    (clk_0),
      .clocks_0_avalon_clocks_slave_readdata_from_sa                          (clocks_0_avalon_clocks_slave_readdata_from_sa),
      .d1_clocks_0_avalon_clocks_slave_end_xfer                               (d1_clocks_0_avalon_clocks_slave_end_xfer),
      .nios_system_clock_9_out_address                                        (nios_system_clock_9_out_address),
      .nios_system_clock_9_out_address_to_slave                               (nios_system_clock_9_out_address_to_slave),
      .nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave           (nios_system_clock_9_out_granted_clocks_0_avalon_clocks_slave),
      .nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave (nios_system_clock_9_out_qualified_request_clocks_0_avalon_clocks_slave),
      .nios_system_clock_9_out_read                                           (nios_system_clock_9_out_read),
      .nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave   (nios_system_clock_9_out_read_data_valid_clocks_0_avalon_clocks_slave),
      .nios_system_clock_9_out_readdata                                       (nios_system_clock_9_out_readdata),
      .nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave          (nios_system_clock_9_out_requests_clocks_0_avalon_clocks_slave),
      .nios_system_clock_9_out_reset_n                                        (nios_system_clock_9_out_reset_n),
      .nios_system_clock_9_out_waitrequest                                    (nios_system_clock_9_out_waitrequest),
      .nios_system_clock_9_out_write                                          (nios_system_clock_9_out_write),
      .nios_system_clock_9_out_writedata                                      (nios_system_clock_9_out_writedata),
      .reset_n                                                                (clk_0_reset_n)
    );

  nios_system_clock_9 the_nios_system_clock_9
    (
      .master_address       (nios_system_clock_9_out_address),
      .master_clk           (clk_0),
      .master_endofpacket   (nios_system_clock_9_out_endofpacket),
      .master_nativeaddress (nios_system_clock_9_out_nativeaddress),
      .master_read          (nios_system_clock_9_out_read),
      .master_readdata      (nios_system_clock_9_out_readdata),
      .master_reset_n       (nios_system_clock_9_out_reset_n),
      .master_waitrequest   (nios_system_clock_9_out_waitrequest),
      .master_write         (nios_system_clock_9_out_write),
      .master_writedata     (nios_system_clock_9_out_writedata),
      .slave_address        (nios_system_clock_9_in_address),
      .slave_clk            (sys_clk),
      .slave_endofpacket    (nios_system_clock_9_in_endofpacket),
      .slave_nativeaddress  (nios_system_clock_9_in_nativeaddress),
      .slave_read           (nios_system_clock_9_in_read),
      .slave_readdata       (nios_system_clock_9_in_readdata),
      .slave_reset_n        (nios_system_clock_9_in_reset_n),
      .slave_waitrequest    (nios_system_clock_9_in_waitrequest),
      .slave_write          (nios_system_clock_9_in_write),
      .slave_writedata      (nios_system_clock_9_in_writedata)
    );

  onchip_memory2_0_s1_arbitrator the_onchip_memory2_0_s1
    (
      .clk                                                                              (sys_clk),
      .cpu_0_data_master_address_to_slave                                               (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                                     (cpu_0_data_master_byteenable),
      .cpu_0_data_master_granted_onchip_memory2_0_s1                                    (cpu_0_data_master_granted_onchip_memory2_0_s1),
      .cpu_0_data_master_latency_counter                                                (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_onchip_memory2_0_s1                          (cpu_0_data_master_qualified_request_onchip_memory2_0_s1),
      .cpu_0_data_master_read                                                           (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_onchip_memory2_0_s1                            (cpu_0_data_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_onchip_memory2_0_s1                                   (cpu_0_data_master_requests_onchip_memory2_0_s1),
      .cpu_0_data_master_write                                                          (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                                      (cpu_0_data_master_writedata),
      .cpu_0_instruction_master_address_to_slave                                        (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_granted_onchip_memory2_0_s1                             (cpu_0_instruction_master_granted_onchip_memory2_0_s1),
      .cpu_0_instruction_master_latency_counter                                         (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1                   (cpu_0_instruction_master_qualified_request_onchip_memory2_0_s1),
      .cpu_0_instruction_master_read                                                    (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1                     (cpu_0_instruction_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_0_instruction_master_requests_onchip_memory2_0_s1                            (cpu_0_instruction_master_requests_onchip_memory2_0_s1),
      .cpu_1_data_master_address_to_slave                                               (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_byteenable                                                     (cpu_1_data_master_byteenable),
      .cpu_1_data_master_granted_onchip_memory2_0_s1                                    (cpu_1_data_master_granted_onchip_memory2_0_s1),
      .cpu_1_data_master_latency_counter                                                (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_onchip_memory2_0_s1                          (cpu_1_data_master_qualified_request_onchip_memory2_0_s1),
      .cpu_1_data_master_read                                                           (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_onchip_memory2_0_s1                            (cpu_1_data_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_onchip_memory2_0_s1                                   (cpu_1_data_master_requests_onchip_memory2_0_s1),
      .cpu_1_data_master_write                                                          (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                                      (cpu_1_data_master_writedata),
      .cpu_1_instruction_master_address_to_slave                                        (cpu_1_instruction_master_address_to_slave),
      .cpu_1_instruction_master_granted_onchip_memory2_0_s1                             (cpu_1_instruction_master_granted_onchip_memory2_0_s1),
      .cpu_1_instruction_master_latency_counter                                         (cpu_1_instruction_master_latency_counter),
      .cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1                   (cpu_1_instruction_master_qualified_request_onchip_memory2_0_s1),
      .cpu_1_instruction_master_read                                                    (cpu_1_instruction_master_read),
      .cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1                     (cpu_1_instruction_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_instruction_master_requests_onchip_memory2_0_s1                            (cpu_1_instruction_master_requests_onchip_memory2_0_s1),
      .cpu_2_data_master_address_to_slave                                               (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_byteenable                                                     (cpu_2_data_master_byteenable),
      .cpu_2_data_master_granted_onchip_memory2_0_s1                                    (cpu_2_data_master_granted_onchip_memory2_0_s1),
      .cpu_2_data_master_latency_counter                                                (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_onchip_memory2_0_s1                          (cpu_2_data_master_qualified_request_onchip_memory2_0_s1),
      .cpu_2_data_master_read                                                           (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_onchip_memory2_0_s1                            (cpu_2_data_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_onchip_memory2_0_s1                                   (cpu_2_data_master_requests_onchip_memory2_0_s1),
      .cpu_2_data_master_write                                                          (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                                      (cpu_2_data_master_writedata),
      .cpu_2_instruction_master_address_to_slave                                        (cpu_2_instruction_master_address_to_slave),
      .cpu_2_instruction_master_granted_onchip_memory2_0_s1                             (cpu_2_instruction_master_granted_onchip_memory2_0_s1),
      .cpu_2_instruction_master_latency_counter                                         (cpu_2_instruction_master_latency_counter),
      .cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1                   (cpu_2_instruction_master_qualified_request_onchip_memory2_0_s1),
      .cpu_2_instruction_master_read                                                    (cpu_2_instruction_master_read),
      .cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1                     (cpu_2_instruction_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_instruction_master_requests_onchip_memory2_0_s1                            (cpu_2_instruction_master_requests_onchip_memory2_0_s1),
      .cpu_3_data_master_address_to_slave                                               (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_byteenable                                                     (cpu_3_data_master_byteenable),
      .cpu_3_data_master_granted_onchip_memory2_0_s1                                    (cpu_3_data_master_granted_onchip_memory2_0_s1),
      .cpu_3_data_master_latency_counter                                                (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_onchip_memory2_0_s1                          (cpu_3_data_master_qualified_request_onchip_memory2_0_s1),
      .cpu_3_data_master_read                                                           (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_onchip_memory2_0_s1                            (cpu_3_data_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_onchip_memory2_0_s1                                   (cpu_3_data_master_requests_onchip_memory2_0_s1),
      .cpu_3_data_master_write                                                          (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                                      (cpu_3_data_master_writedata),
      .cpu_3_instruction_master_address_to_slave                                        (cpu_3_instruction_master_address_to_slave),
      .cpu_3_instruction_master_granted_onchip_memory2_0_s1                             (cpu_3_instruction_master_granted_onchip_memory2_0_s1),
      .cpu_3_instruction_master_latency_counter                                         (cpu_3_instruction_master_latency_counter),
      .cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1                   (cpu_3_instruction_master_qualified_request_onchip_memory2_0_s1),
      .cpu_3_instruction_master_read                                                    (cpu_3_instruction_master_read),
      .cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1                     (cpu_3_instruction_master_read_data_valid_onchip_memory2_0_s1),
      .cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_instruction_master_requests_onchip_memory2_0_s1                            (cpu_3_instruction_master_requests_onchip_memory2_0_s1),
      .d1_onchip_memory2_0_s1_end_xfer                                                  (d1_onchip_memory2_0_s1_end_xfer),
      .onchip_memory2_0_s1_address                                                      (onchip_memory2_0_s1_address),
      .onchip_memory2_0_s1_byteenable                                                   (onchip_memory2_0_s1_byteenable),
      .onchip_memory2_0_s1_chipselect                                                   (onchip_memory2_0_s1_chipselect),
      .onchip_memory2_0_s1_clken                                                        (onchip_memory2_0_s1_clken),
      .onchip_memory2_0_s1_readdata                                                     (onchip_memory2_0_s1_readdata),
      .onchip_memory2_0_s1_readdata_from_sa                                             (onchip_memory2_0_s1_readdata_from_sa),
      .onchip_memory2_0_s1_reset                                                        (onchip_memory2_0_s1_reset),
      .onchip_memory2_0_s1_write                                                        (onchip_memory2_0_s1_write),
      .onchip_memory2_0_s1_writedata                                                    (onchip_memory2_0_s1_writedata),
      .reset_n                                                                          (sys_clk_reset_n)
    );

  onchip_memory2_0 the_onchip_memory2_0
    (
      .address    (onchip_memory2_0_s1_address),
      .byteenable (onchip_memory2_0_s1_byteenable),
      .chipselect (onchip_memory2_0_s1_chipselect),
      .clk        (sys_clk),
      .clken      (onchip_memory2_0_s1_clken),
      .readdata   (onchip_memory2_0_s1_readdata),
      .reset      (onchip_memory2_0_s1_reset),
      .write      (onchip_memory2_0_s1_write),
      .writedata  (onchip_memory2_0_s1_writedata)
    );

  onchip_memory2_1_s1_arbitrator the_onchip_memory2_1_s1
    (
      .clk                                                                              (sys_clk),
      .cpu_0_data_master_address_to_slave                                               (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                                     (cpu_0_data_master_byteenable),
      .cpu_0_data_master_granted_onchip_memory2_1_s1                                    (cpu_0_data_master_granted_onchip_memory2_1_s1),
      .cpu_0_data_master_latency_counter                                                (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_onchip_memory2_1_s1                          (cpu_0_data_master_qualified_request_onchip_memory2_1_s1),
      .cpu_0_data_master_read                                                           (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_onchip_memory2_1_s1                            (cpu_0_data_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_onchip_memory2_1_s1                                   (cpu_0_data_master_requests_onchip_memory2_1_s1),
      .cpu_0_data_master_write                                                          (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                                      (cpu_0_data_master_writedata),
      .cpu_0_instruction_master_address_to_slave                                        (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_granted_onchip_memory2_1_s1                             (cpu_0_instruction_master_granted_onchip_memory2_1_s1),
      .cpu_0_instruction_master_latency_counter                                         (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1                   (cpu_0_instruction_master_qualified_request_onchip_memory2_1_s1),
      .cpu_0_instruction_master_read                                                    (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1                     (cpu_0_instruction_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_0_instruction_master_requests_onchip_memory2_1_s1                            (cpu_0_instruction_master_requests_onchip_memory2_1_s1),
      .cpu_1_data_master_address_to_slave                                               (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_byteenable                                                     (cpu_1_data_master_byteenable),
      .cpu_1_data_master_granted_onchip_memory2_1_s1                                    (cpu_1_data_master_granted_onchip_memory2_1_s1),
      .cpu_1_data_master_latency_counter                                                (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_onchip_memory2_1_s1                          (cpu_1_data_master_qualified_request_onchip_memory2_1_s1),
      .cpu_1_data_master_read                                                           (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_onchip_memory2_1_s1                            (cpu_1_data_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_onchip_memory2_1_s1                                   (cpu_1_data_master_requests_onchip_memory2_1_s1),
      .cpu_1_data_master_write                                                          (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                                      (cpu_1_data_master_writedata),
      .cpu_1_instruction_master_address_to_slave                                        (cpu_1_instruction_master_address_to_slave),
      .cpu_1_instruction_master_granted_onchip_memory2_1_s1                             (cpu_1_instruction_master_granted_onchip_memory2_1_s1),
      .cpu_1_instruction_master_latency_counter                                         (cpu_1_instruction_master_latency_counter),
      .cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1                   (cpu_1_instruction_master_qualified_request_onchip_memory2_1_s1),
      .cpu_1_instruction_master_read                                                    (cpu_1_instruction_master_read),
      .cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1                     (cpu_1_instruction_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_instruction_master_requests_onchip_memory2_1_s1                            (cpu_1_instruction_master_requests_onchip_memory2_1_s1),
      .cpu_2_data_master_address_to_slave                                               (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_byteenable                                                     (cpu_2_data_master_byteenable),
      .cpu_2_data_master_granted_onchip_memory2_1_s1                                    (cpu_2_data_master_granted_onchip_memory2_1_s1),
      .cpu_2_data_master_latency_counter                                                (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_onchip_memory2_1_s1                          (cpu_2_data_master_qualified_request_onchip_memory2_1_s1),
      .cpu_2_data_master_read                                                           (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_onchip_memory2_1_s1                            (cpu_2_data_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_onchip_memory2_1_s1                                   (cpu_2_data_master_requests_onchip_memory2_1_s1),
      .cpu_2_data_master_write                                                          (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                                      (cpu_2_data_master_writedata),
      .cpu_2_instruction_master_address_to_slave                                        (cpu_2_instruction_master_address_to_slave),
      .cpu_2_instruction_master_granted_onchip_memory2_1_s1                             (cpu_2_instruction_master_granted_onchip_memory2_1_s1),
      .cpu_2_instruction_master_latency_counter                                         (cpu_2_instruction_master_latency_counter),
      .cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1                   (cpu_2_instruction_master_qualified_request_onchip_memory2_1_s1),
      .cpu_2_instruction_master_read                                                    (cpu_2_instruction_master_read),
      .cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1                     (cpu_2_instruction_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_instruction_master_requests_onchip_memory2_1_s1                            (cpu_2_instruction_master_requests_onchip_memory2_1_s1),
      .cpu_3_data_master_address_to_slave                                               (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_byteenable                                                     (cpu_3_data_master_byteenable),
      .cpu_3_data_master_granted_onchip_memory2_1_s1                                    (cpu_3_data_master_granted_onchip_memory2_1_s1),
      .cpu_3_data_master_latency_counter                                                (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_onchip_memory2_1_s1                          (cpu_3_data_master_qualified_request_onchip_memory2_1_s1),
      .cpu_3_data_master_read                                                           (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_onchip_memory2_1_s1                            (cpu_3_data_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_onchip_memory2_1_s1                                   (cpu_3_data_master_requests_onchip_memory2_1_s1),
      .cpu_3_data_master_write                                                          (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                                      (cpu_3_data_master_writedata),
      .cpu_3_instruction_master_address_to_slave                                        (cpu_3_instruction_master_address_to_slave),
      .cpu_3_instruction_master_granted_onchip_memory2_1_s1                             (cpu_3_instruction_master_granted_onchip_memory2_1_s1),
      .cpu_3_instruction_master_latency_counter                                         (cpu_3_instruction_master_latency_counter),
      .cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1                   (cpu_3_instruction_master_qualified_request_onchip_memory2_1_s1),
      .cpu_3_instruction_master_read                                                    (cpu_3_instruction_master_read),
      .cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1                     (cpu_3_instruction_master_read_data_valid_onchip_memory2_1_s1),
      .cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_instruction_master_requests_onchip_memory2_1_s1                            (cpu_3_instruction_master_requests_onchip_memory2_1_s1),
      .d1_onchip_memory2_1_s1_end_xfer                                                  (d1_onchip_memory2_1_s1_end_xfer),
      .onchip_memory2_1_s1_address                                                      (onchip_memory2_1_s1_address),
      .onchip_memory2_1_s1_byteenable                                                   (onchip_memory2_1_s1_byteenable),
      .onchip_memory2_1_s1_chipselect                                                   (onchip_memory2_1_s1_chipselect),
      .onchip_memory2_1_s1_clken                                                        (onchip_memory2_1_s1_clken),
      .onchip_memory2_1_s1_readdata                                                     (onchip_memory2_1_s1_readdata),
      .onchip_memory2_1_s1_readdata_from_sa                                             (onchip_memory2_1_s1_readdata_from_sa),
      .onchip_memory2_1_s1_reset                                                        (onchip_memory2_1_s1_reset),
      .onchip_memory2_1_s1_write                                                        (onchip_memory2_1_s1_write),
      .onchip_memory2_1_s1_writedata                                                    (onchip_memory2_1_s1_writedata),
      .reset_n                                                                          (sys_clk_reset_n)
    );

  onchip_memory2_1 the_onchip_memory2_1
    (
      .address    (onchip_memory2_1_s1_address),
      .byteenable (onchip_memory2_1_s1_byteenable),
      .chipselect (onchip_memory2_1_s1_chipselect),
      .clk        (sys_clk),
      .clken      (onchip_memory2_1_s1_clken),
      .readdata   (onchip_memory2_1_s1_readdata),
      .reset      (onchip_memory2_1_s1_reset),
      .write      (onchip_memory2_1_s1_write),
      .writedata  (onchip_memory2_1_s1_writedata)
    );

  onchip_memory2_2_s1_arbitrator the_onchip_memory2_2_s1
    (
      .clk                                                                              (sys_clk),
      .cpu_0_data_master_address_to_slave                                               (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                                     (cpu_0_data_master_byteenable),
      .cpu_0_data_master_granted_onchip_memory2_2_s1                                    (cpu_0_data_master_granted_onchip_memory2_2_s1),
      .cpu_0_data_master_latency_counter                                                (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_onchip_memory2_2_s1                          (cpu_0_data_master_qualified_request_onchip_memory2_2_s1),
      .cpu_0_data_master_read                                                           (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_onchip_memory2_2_s1                            (cpu_0_data_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_onchip_memory2_2_s1                                   (cpu_0_data_master_requests_onchip_memory2_2_s1),
      .cpu_0_data_master_write                                                          (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                                      (cpu_0_data_master_writedata),
      .cpu_0_instruction_master_address_to_slave                                        (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_granted_onchip_memory2_2_s1                             (cpu_0_instruction_master_granted_onchip_memory2_2_s1),
      .cpu_0_instruction_master_latency_counter                                         (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1                   (cpu_0_instruction_master_qualified_request_onchip_memory2_2_s1),
      .cpu_0_instruction_master_read                                                    (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1                     (cpu_0_instruction_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_0_instruction_master_requests_onchip_memory2_2_s1                            (cpu_0_instruction_master_requests_onchip_memory2_2_s1),
      .cpu_1_data_master_address_to_slave                                               (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_byteenable                                                     (cpu_1_data_master_byteenable),
      .cpu_1_data_master_granted_onchip_memory2_2_s1                                    (cpu_1_data_master_granted_onchip_memory2_2_s1),
      .cpu_1_data_master_latency_counter                                                (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_onchip_memory2_2_s1                          (cpu_1_data_master_qualified_request_onchip_memory2_2_s1),
      .cpu_1_data_master_read                                                           (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_onchip_memory2_2_s1                            (cpu_1_data_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_onchip_memory2_2_s1                                   (cpu_1_data_master_requests_onchip_memory2_2_s1),
      .cpu_1_data_master_write                                                          (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                                      (cpu_1_data_master_writedata),
      .cpu_1_instruction_master_address_to_slave                                        (cpu_1_instruction_master_address_to_slave),
      .cpu_1_instruction_master_granted_onchip_memory2_2_s1                             (cpu_1_instruction_master_granted_onchip_memory2_2_s1),
      .cpu_1_instruction_master_latency_counter                                         (cpu_1_instruction_master_latency_counter),
      .cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1                   (cpu_1_instruction_master_qualified_request_onchip_memory2_2_s1),
      .cpu_1_instruction_master_read                                                    (cpu_1_instruction_master_read),
      .cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1                     (cpu_1_instruction_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_instruction_master_requests_onchip_memory2_2_s1                            (cpu_1_instruction_master_requests_onchip_memory2_2_s1),
      .cpu_2_data_master_address_to_slave                                               (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_byteenable                                                     (cpu_2_data_master_byteenable),
      .cpu_2_data_master_granted_onchip_memory2_2_s1                                    (cpu_2_data_master_granted_onchip_memory2_2_s1),
      .cpu_2_data_master_latency_counter                                                (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_onchip_memory2_2_s1                          (cpu_2_data_master_qualified_request_onchip_memory2_2_s1),
      .cpu_2_data_master_read                                                           (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_onchip_memory2_2_s1                            (cpu_2_data_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_onchip_memory2_2_s1                                   (cpu_2_data_master_requests_onchip_memory2_2_s1),
      .cpu_2_data_master_write                                                          (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                                      (cpu_2_data_master_writedata),
      .cpu_2_instruction_master_address_to_slave                                        (cpu_2_instruction_master_address_to_slave),
      .cpu_2_instruction_master_granted_onchip_memory2_2_s1                             (cpu_2_instruction_master_granted_onchip_memory2_2_s1),
      .cpu_2_instruction_master_latency_counter                                         (cpu_2_instruction_master_latency_counter),
      .cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1                   (cpu_2_instruction_master_qualified_request_onchip_memory2_2_s1),
      .cpu_2_instruction_master_read                                                    (cpu_2_instruction_master_read),
      .cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1                     (cpu_2_instruction_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_instruction_master_requests_onchip_memory2_2_s1                            (cpu_2_instruction_master_requests_onchip_memory2_2_s1),
      .cpu_3_data_master_address_to_slave                                               (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_byteenable                                                     (cpu_3_data_master_byteenable),
      .cpu_3_data_master_granted_onchip_memory2_2_s1                                    (cpu_3_data_master_granted_onchip_memory2_2_s1),
      .cpu_3_data_master_latency_counter                                                (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_onchip_memory2_2_s1                          (cpu_3_data_master_qualified_request_onchip_memory2_2_s1),
      .cpu_3_data_master_read                                                           (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_onchip_memory2_2_s1                            (cpu_3_data_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_onchip_memory2_2_s1                                   (cpu_3_data_master_requests_onchip_memory2_2_s1),
      .cpu_3_data_master_write                                                          (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                                      (cpu_3_data_master_writedata),
      .cpu_3_instruction_master_address_to_slave                                        (cpu_3_instruction_master_address_to_slave),
      .cpu_3_instruction_master_granted_onchip_memory2_2_s1                             (cpu_3_instruction_master_granted_onchip_memory2_2_s1),
      .cpu_3_instruction_master_latency_counter                                         (cpu_3_instruction_master_latency_counter),
      .cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1                   (cpu_3_instruction_master_qualified_request_onchip_memory2_2_s1),
      .cpu_3_instruction_master_read                                                    (cpu_3_instruction_master_read),
      .cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1                     (cpu_3_instruction_master_read_data_valid_onchip_memory2_2_s1),
      .cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_instruction_master_requests_onchip_memory2_2_s1                            (cpu_3_instruction_master_requests_onchip_memory2_2_s1),
      .d1_onchip_memory2_2_s1_end_xfer                                                  (d1_onchip_memory2_2_s1_end_xfer),
      .onchip_memory2_2_s1_address                                                      (onchip_memory2_2_s1_address),
      .onchip_memory2_2_s1_byteenable                                                   (onchip_memory2_2_s1_byteenable),
      .onchip_memory2_2_s1_chipselect                                                   (onchip_memory2_2_s1_chipselect),
      .onchip_memory2_2_s1_clken                                                        (onchip_memory2_2_s1_clken),
      .onchip_memory2_2_s1_readdata                                                     (onchip_memory2_2_s1_readdata),
      .onchip_memory2_2_s1_readdata_from_sa                                             (onchip_memory2_2_s1_readdata_from_sa),
      .onchip_memory2_2_s1_reset                                                        (onchip_memory2_2_s1_reset),
      .onchip_memory2_2_s1_write                                                        (onchip_memory2_2_s1_write),
      .onchip_memory2_2_s1_writedata                                                    (onchip_memory2_2_s1_writedata),
      .reset_n                                                                          (sys_clk_reset_n)
    );

  onchip_memory2_2 the_onchip_memory2_2
    (
      .address    (onchip_memory2_2_s1_address),
      .byteenable (onchip_memory2_2_s1_byteenable),
      .chipselect (onchip_memory2_2_s1_chipselect),
      .clk        (sys_clk),
      .clken      (onchip_memory2_2_s1_clken),
      .readdata   (onchip_memory2_2_s1_readdata),
      .reset      (onchip_memory2_2_s1_reset),
      .write      (onchip_memory2_2_s1_write),
      .writedata  (onchip_memory2_2_s1_writedata)
    );

  onchip_memory2_3_s1_arbitrator the_onchip_memory2_3_s1
    (
      .clk                                                                              (sys_clk),
      .cpu_0_data_master_address_to_slave                                               (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                                     (cpu_0_data_master_byteenable),
      .cpu_0_data_master_granted_onchip_memory2_3_s1                                    (cpu_0_data_master_granted_onchip_memory2_3_s1),
      .cpu_0_data_master_latency_counter                                                (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_onchip_memory2_3_s1                          (cpu_0_data_master_qualified_request_onchip_memory2_3_s1),
      .cpu_0_data_master_read                                                           (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_onchip_memory2_3_s1                            (cpu_0_data_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_onchip_memory2_3_s1                                   (cpu_0_data_master_requests_onchip_memory2_3_s1),
      .cpu_0_data_master_write                                                          (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                                      (cpu_0_data_master_writedata),
      .cpu_0_instruction_master_address_to_slave                                        (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_granted_onchip_memory2_3_s1                             (cpu_0_instruction_master_granted_onchip_memory2_3_s1),
      .cpu_0_instruction_master_latency_counter                                         (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1                   (cpu_0_instruction_master_qualified_request_onchip_memory2_3_s1),
      .cpu_0_instruction_master_read                                                    (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1                     (cpu_0_instruction_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_0_instruction_master_requests_onchip_memory2_3_s1                            (cpu_0_instruction_master_requests_onchip_memory2_3_s1),
      .cpu_1_data_master_address_to_slave                                               (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_byteenable                                                     (cpu_1_data_master_byteenable),
      .cpu_1_data_master_granted_onchip_memory2_3_s1                                    (cpu_1_data_master_granted_onchip_memory2_3_s1),
      .cpu_1_data_master_latency_counter                                                (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_onchip_memory2_3_s1                          (cpu_1_data_master_qualified_request_onchip_memory2_3_s1),
      .cpu_1_data_master_read                                                           (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_onchip_memory2_3_s1                            (cpu_1_data_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_onchip_memory2_3_s1                                   (cpu_1_data_master_requests_onchip_memory2_3_s1),
      .cpu_1_data_master_write                                                          (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                                      (cpu_1_data_master_writedata),
      .cpu_1_instruction_master_address_to_slave                                        (cpu_1_instruction_master_address_to_slave),
      .cpu_1_instruction_master_granted_onchip_memory2_3_s1                             (cpu_1_instruction_master_granted_onchip_memory2_3_s1),
      .cpu_1_instruction_master_latency_counter                                         (cpu_1_instruction_master_latency_counter),
      .cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1                   (cpu_1_instruction_master_qualified_request_onchip_memory2_3_s1),
      .cpu_1_instruction_master_read                                                    (cpu_1_instruction_master_read),
      .cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1                     (cpu_1_instruction_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_instruction_master_requests_onchip_memory2_3_s1                            (cpu_1_instruction_master_requests_onchip_memory2_3_s1),
      .cpu_2_data_master_address_to_slave                                               (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_byteenable                                                     (cpu_2_data_master_byteenable),
      .cpu_2_data_master_granted_onchip_memory2_3_s1                                    (cpu_2_data_master_granted_onchip_memory2_3_s1),
      .cpu_2_data_master_latency_counter                                                (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_onchip_memory2_3_s1                          (cpu_2_data_master_qualified_request_onchip_memory2_3_s1),
      .cpu_2_data_master_read                                                           (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_onchip_memory2_3_s1                            (cpu_2_data_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_onchip_memory2_3_s1                                   (cpu_2_data_master_requests_onchip_memory2_3_s1),
      .cpu_2_data_master_write                                                          (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                                      (cpu_2_data_master_writedata),
      .cpu_2_instruction_master_address_to_slave                                        (cpu_2_instruction_master_address_to_slave),
      .cpu_2_instruction_master_granted_onchip_memory2_3_s1                             (cpu_2_instruction_master_granted_onchip_memory2_3_s1),
      .cpu_2_instruction_master_latency_counter                                         (cpu_2_instruction_master_latency_counter),
      .cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1                   (cpu_2_instruction_master_qualified_request_onchip_memory2_3_s1),
      .cpu_2_instruction_master_read                                                    (cpu_2_instruction_master_read),
      .cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1                     (cpu_2_instruction_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_instruction_master_requests_onchip_memory2_3_s1                            (cpu_2_instruction_master_requests_onchip_memory2_3_s1),
      .cpu_3_data_master_address_to_slave                                               (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_byteenable                                                     (cpu_3_data_master_byteenable),
      .cpu_3_data_master_granted_onchip_memory2_3_s1                                    (cpu_3_data_master_granted_onchip_memory2_3_s1),
      .cpu_3_data_master_latency_counter                                                (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_onchip_memory2_3_s1                          (cpu_3_data_master_qualified_request_onchip_memory2_3_s1),
      .cpu_3_data_master_read                                                           (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_onchip_memory2_3_s1                            (cpu_3_data_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register        (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_onchip_memory2_3_s1                                   (cpu_3_data_master_requests_onchip_memory2_3_s1),
      .cpu_3_data_master_write                                                          (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                                      (cpu_3_data_master_writedata),
      .cpu_3_instruction_master_address_to_slave                                        (cpu_3_instruction_master_address_to_slave),
      .cpu_3_instruction_master_granted_onchip_memory2_3_s1                             (cpu_3_instruction_master_granted_onchip_memory2_3_s1),
      .cpu_3_instruction_master_latency_counter                                         (cpu_3_instruction_master_latency_counter),
      .cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1                   (cpu_3_instruction_master_qualified_request_onchip_memory2_3_s1),
      .cpu_3_instruction_master_read                                                    (cpu_3_instruction_master_read),
      .cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1                     (cpu_3_instruction_master_read_data_valid_onchip_memory2_3_s1),
      .cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_instruction_master_requests_onchip_memory2_3_s1                            (cpu_3_instruction_master_requests_onchip_memory2_3_s1),
      .d1_onchip_memory2_3_s1_end_xfer                                                  (d1_onchip_memory2_3_s1_end_xfer),
      .onchip_memory2_3_s1_address                                                      (onchip_memory2_3_s1_address),
      .onchip_memory2_3_s1_byteenable                                                   (onchip_memory2_3_s1_byteenable),
      .onchip_memory2_3_s1_chipselect                                                   (onchip_memory2_3_s1_chipselect),
      .onchip_memory2_3_s1_clken                                                        (onchip_memory2_3_s1_clken),
      .onchip_memory2_3_s1_readdata                                                     (onchip_memory2_3_s1_readdata),
      .onchip_memory2_3_s1_readdata_from_sa                                             (onchip_memory2_3_s1_readdata_from_sa),
      .onchip_memory2_3_s1_reset                                                        (onchip_memory2_3_s1_reset),
      .onchip_memory2_3_s1_write                                                        (onchip_memory2_3_s1_write),
      .onchip_memory2_3_s1_writedata                                                    (onchip_memory2_3_s1_writedata),
      .reset_n                                                                          (sys_clk_reset_n)
    );

  onchip_memory2_3 the_onchip_memory2_3
    (
      .address    (onchip_memory2_3_s1_address),
      .byteenable (onchip_memory2_3_s1_byteenable),
      .chipselect (onchip_memory2_3_s1_chipselect),
      .clk        (sys_clk),
      .clken      (onchip_memory2_3_s1_clken),
      .readdata   (onchip_memory2_3_s1_readdata),
      .reset      (onchip_memory2_3_s1_reset),
      .write      (onchip_memory2_3_s1_write),
      .writedata  (onchip_memory2_3_s1_writedata)
    );

  performance_counter_0_control_slave_arbitrator the_performance_counter_0_control_slave
    (
      .clk                                                                       (sys_clk),
      .cpu_0_data_master_address_to_slave                                        (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_performance_counter_0_control_slave             (cpu_0_data_master_granted_performance_counter_0_control_slave),
      .cpu_0_data_master_latency_counter                                         (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_performance_counter_0_control_slave   (cpu_0_data_master_qualified_request_performance_counter_0_control_slave),
      .cpu_0_data_master_read                                                    (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_performance_counter_0_control_slave     (cpu_0_data_master_read_data_valid_performance_counter_0_control_slave),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_performance_counter_0_control_slave            (cpu_0_data_master_requests_performance_counter_0_control_slave),
      .cpu_0_data_master_write                                                   (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                               (cpu_0_data_master_writedata),
      .cpu_1_data_master_address_to_slave                                        (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_granted_performance_counter_0_control_slave             (cpu_1_data_master_granted_performance_counter_0_control_slave),
      .cpu_1_data_master_latency_counter                                         (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_performance_counter_0_control_slave   (cpu_1_data_master_qualified_request_performance_counter_0_control_slave),
      .cpu_1_data_master_read                                                    (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_performance_counter_0_control_slave     (cpu_1_data_master_read_data_valid_performance_counter_0_control_slave),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_performance_counter_0_control_slave            (cpu_1_data_master_requests_performance_counter_0_control_slave),
      .cpu_1_data_master_write                                                   (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                               (cpu_1_data_master_writedata),
      .cpu_2_data_master_address_to_slave                                        (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_granted_performance_counter_0_control_slave             (cpu_2_data_master_granted_performance_counter_0_control_slave),
      .cpu_2_data_master_latency_counter                                         (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_performance_counter_0_control_slave   (cpu_2_data_master_qualified_request_performance_counter_0_control_slave),
      .cpu_2_data_master_read                                                    (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_performance_counter_0_control_slave     (cpu_2_data_master_read_data_valid_performance_counter_0_control_slave),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_performance_counter_0_control_slave            (cpu_2_data_master_requests_performance_counter_0_control_slave),
      .cpu_2_data_master_write                                                   (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                               (cpu_2_data_master_writedata),
      .cpu_3_data_master_address_to_slave                                        (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_granted_performance_counter_0_control_slave             (cpu_3_data_master_granted_performance_counter_0_control_slave),
      .cpu_3_data_master_latency_counter                                         (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_performance_counter_0_control_slave   (cpu_3_data_master_qualified_request_performance_counter_0_control_slave),
      .cpu_3_data_master_read                                                    (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_performance_counter_0_control_slave     (cpu_3_data_master_read_data_valid_performance_counter_0_control_slave),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_performance_counter_0_control_slave            (cpu_3_data_master_requests_performance_counter_0_control_slave),
      .cpu_3_data_master_write                                                   (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                               (cpu_3_data_master_writedata),
      .d1_performance_counter_0_control_slave_end_xfer                           (d1_performance_counter_0_control_slave_end_xfer),
      .performance_counter_0_control_slave_address                               (performance_counter_0_control_slave_address),
      .performance_counter_0_control_slave_begintransfer                         (performance_counter_0_control_slave_begintransfer),
      .performance_counter_0_control_slave_readdata                              (performance_counter_0_control_slave_readdata),
      .performance_counter_0_control_slave_readdata_from_sa                      (performance_counter_0_control_slave_readdata_from_sa),
      .performance_counter_0_control_slave_reset_n                               (performance_counter_0_control_slave_reset_n),
      .performance_counter_0_control_slave_write                                 (performance_counter_0_control_slave_write),
      .performance_counter_0_control_slave_writedata                             (performance_counter_0_control_slave_writedata),
      .reset_n                                                                   (sys_clk_reset_n)
    );

  performance_counter_0 the_performance_counter_0
    (
      .address       (performance_counter_0_control_slave_address),
      .begintransfer (performance_counter_0_control_slave_begintransfer),
      .clk           (sys_clk),
      .readdata      (performance_counter_0_control_slave_readdata),
      .reset_n       (performance_counter_0_control_slave_reset_n),
      .write         (performance_counter_0_control_slave_write),
      .writedata     (performance_counter_0_control_slave_writedata)
    );

  sdram_0_s1_arbitrator the_sdram_0_s1
    (
      .clk                                                               (sdram_clk),
      .d1_sdram_0_s1_end_xfer                                            (d1_sdram_0_s1_end_xfer),
      .nios_system_clock_0_out_address_to_slave                          (nios_system_clock_0_out_address_to_slave),
      .nios_system_clock_0_out_byteenable                                (nios_system_clock_0_out_byteenable),
      .nios_system_clock_0_out_granted_sdram_0_s1                        (nios_system_clock_0_out_granted_sdram_0_s1),
      .nios_system_clock_0_out_qualified_request_sdram_0_s1              (nios_system_clock_0_out_qualified_request_sdram_0_s1),
      .nios_system_clock_0_out_read                                      (nios_system_clock_0_out_read),
      .nios_system_clock_0_out_read_data_valid_sdram_0_s1                (nios_system_clock_0_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_0_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_0_out_requests_sdram_0_s1                       (nios_system_clock_0_out_requests_sdram_0_s1),
      .nios_system_clock_0_out_write                                     (nios_system_clock_0_out_write),
      .nios_system_clock_0_out_writedata                                 (nios_system_clock_0_out_writedata),
      .nios_system_clock_1_out_address_to_slave                          (nios_system_clock_1_out_address_to_slave),
      .nios_system_clock_1_out_byteenable                                (nios_system_clock_1_out_byteenable),
      .nios_system_clock_1_out_granted_sdram_0_s1                        (nios_system_clock_1_out_granted_sdram_0_s1),
      .nios_system_clock_1_out_qualified_request_sdram_0_s1              (nios_system_clock_1_out_qualified_request_sdram_0_s1),
      .nios_system_clock_1_out_read                                      (nios_system_clock_1_out_read),
      .nios_system_clock_1_out_read_data_valid_sdram_0_s1                (nios_system_clock_1_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_1_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_1_out_requests_sdram_0_s1                       (nios_system_clock_1_out_requests_sdram_0_s1),
      .nios_system_clock_1_out_write                                     (nios_system_clock_1_out_write),
      .nios_system_clock_1_out_writedata                                 (nios_system_clock_1_out_writedata),
      .nios_system_clock_2_out_address_to_slave                          (nios_system_clock_2_out_address_to_slave),
      .nios_system_clock_2_out_byteenable                                (nios_system_clock_2_out_byteenable),
      .nios_system_clock_2_out_granted_sdram_0_s1                        (nios_system_clock_2_out_granted_sdram_0_s1),
      .nios_system_clock_2_out_qualified_request_sdram_0_s1              (nios_system_clock_2_out_qualified_request_sdram_0_s1),
      .nios_system_clock_2_out_read                                      (nios_system_clock_2_out_read),
      .nios_system_clock_2_out_read_data_valid_sdram_0_s1                (nios_system_clock_2_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_2_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_2_out_requests_sdram_0_s1                       (nios_system_clock_2_out_requests_sdram_0_s1),
      .nios_system_clock_2_out_write                                     (nios_system_clock_2_out_write),
      .nios_system_clock_2_out_writedata                                 (nios_system_clock_2_out_writedata),
      .nios_system_clock_3_out_address_to_slave                          (nios_system_clock_3_out_address_to_slave),
      .nios_system_clock_3_out_byteenable                                (nios_system_clock_3_out_byteenable),
      .nios_system_clock_3_out_granted_sdram_0_s1                        (nios_system_clock_3_out_granted_sdram_0_s1),
      .nios_system_clock_3_out_qualified_request_sdram_0_s1              (nios_system_clock_3_out_qualified_request_sdram_0_s1),
      .nios_system_clock_3_out_read                                      (nios_system_clock_3_out_read),
      .nios_system_clock_3_out_read_data_valid_sdram_0_s1                (nios_system_clock_3_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_3_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_3_out_requests_sdram_0_s1                       (nios_system_clock_3_out_requests_sdram_0_s1),
      .nios_system_clock_3_out_write                                     (nios_system_clock_3_out_write),
      .nios_system_clock_3_out_writedata                                 (nios_system_clock_3_out_writedata),
      .nios_system_clock_4_out_address_to_slave                          (nios_system_clock_4_out_address_to_slave),
      .nios_system_clock_4_out_byteenable                                (nios_system_clock_4_out_byteenable),
      .nios_system_clock_4_out_granted_sdram_0_s1                        (nios_system_clock_4_out_granted_sdram_0_s1),
      .nios_system_clock_4_out_qualified_request_sdram_0_s1              (nios_system_clock_4_out_qualified_request_sdram_0_s1),
      .nios_system_clock_4_out_read                                      (nios_system_clock_4_out_read),
      .nios_system_clock_4_out_read_data_valid_sdram_0_s1                (nios_system_clock_4_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_4_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_4_out_requests_sdram_0_s1                       (nios_system_clock_4_out_requests_sdram_0_s1),
      .nios_system_clock_4_out_write                                     (nios_system_clock_4_out_write),
      .nios_system_clock_4_out_writedata                                 (nios_system_clock_4_out_writedata),
      .nios_system_clock_5_out_address_to_slave                          (nios_system_clock_5_out_address_to_slave),
      .nios_system_clock_5_out_byteenable                                (nios_system_clock_5_out_byteenable),
      .nios_system_clock_5_out_granted_sdram_0_s1                        (nios_system_clock_5_out_granted_sdram_0_s1),
      .nios_system_clock_5_out_qualified_request_sdram_0_s1              (nios_system_clock_5_out_qualified_request_sdram_0_s1),
      .nios_system_clock_5_out_read                                      (nios_system_clock_5_out_read),
      .nios_system_clock_5_out_read_data_valid_sdram_0_s1                (nios_system_clock_5_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_5_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_5_out_requests_sdram_0_s1                       (nios_system_clock_5_out_requests_sdram_0_s1),
      .nios_system_clock_5_out_write                                     (nios_system_clock_5_out_write),
      .nios_system_clock_5_out_writedata                                 (nios_system_clock_5_out_writedata),
      .nios_system_clock_6_out_address_to_slave                          (nios_system_clock_6_out_address_to_slave),
      .nios_system_clock_6_out_byteenable                                (nios_system_clock_6_out_byteenable),
      .nios_system_clock_6_out_granted_sdram_0_s1                        (nios_system_clock_6_out_granted_sdram_0_s1),
      .nios_system_clock_6_out_qualified_request_sdram_0_s1              (nios_system_clock_6_out_qualified_request_sdram_0_s1),
      .nios_system_clock_6_out_read                                      (nios_system_clock_6_out_read),
      .nios_system_clock_6_out_read_data_valid_sdram_0_s1                (nios_system_clock_6_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_6_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_6_out_requests_sdram_0_s1                       (nios_system_clock_6_out_requests_sdram_0_s1),
      .nios_system_clock_6_out_write                                     (nios_system_clock_6_out_write),
      .nios_system_clock_6_out_writedata                                 (nios_system_clock_6_out_writedata),
      .nios_system_clock_7_out_address_to_slave                          (nios_system_clock_7_out_address_to_slave),
      .nios_system_clock_7_out_byteenable                                (nios_system_clock_7_out_byteenable),
      .nios_system_clock_7_out_granted_sdram_0_s1                        (nios_system_clock_7_out_granted_sdram_0_s1),
      .nios_system_clock_7_out_qualified_request_sdram_0_s1              (nios_system_clock_7_out_qualified_request_sdram_0_s1),
      .nios_system_clock_7_out_read                                      (nios_system_clock_7_out_read),
      .nios_system_clock_7_out_read_data_valid_sdram_0_s1                (nios_system_clock_7_out_read_data_valid_sdram_0_s1),
      .nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register (nios_system_clock_7_out_read_data_valid_sdram_0_s1_shift_register),
      .nios_system_clock_7_out_requests_sdram_0_s1                       (nios_system_clock_7_out_requests_sdram_0_s1),
      .nios_system_clock_7_out_write                                     (nios_system_clock_7_out_write),
      .nios_system_clock_7_out_writedata                                 (nios_system_clock_7_out_writedata),
      .reset_n                                                           (sdram_clk_reset_n),
      .sdram_0_s1_address                                                (sdram_0_s1_address),
      .sdram_0_s1_byteenable_n                                           (sdram_0_s1_byteenable_n),
      .sdram_0_s1_chipselect                                             (sdram_0_s1_chipselect),
      .sdram_0_s1_read_n                                                 (sdram_0_s1_read_n),
      .sdram_0_s1_readdata                                               (sdram_0_s1_readdata),
      .sdram_0_s1_readdata_from_sa                                       (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_readdatavalid                                          (sdram_0_s1_readdatavalid),
      .sdram_0_s1_reset_n                                                (sdram_0_s1_reset_n),
      .sdram_0_s1_waitrequest                                            (sdram_0_s1_waitrequest),
      .sdram_0_s1_waitrequest_from_sa                                    (sdram_0_s1_waitrequest_from_sa),
      .sdram_0_s1_write_n                                                (sdram_0_s1_write_n),
      .sdram_0_s1_writedata                                              (sdram_0_s1_writedata)
    );

  sdram_0 the_sdram_0
    (
      .az_addr        (sdram_0_s1_address),
      .az_be_n        (sdram_0_s1_byteenable_n),
      .az_cs          (sdram_0_s1_chipselect),
      .az_data        (sdram_0_s1_writedata),
      .az_rd_n        (sdram_0_s1_read_n),
      .az_wr_n        (sdram_0_s1_write_n),
      .clk            (sdram_clk),
      .reset_n        (sdram_0_s1_reset_n),
      .za_data        (sdram_0_s1_readdata),
      .za_valid       (sdram_0_s1_readdatavalid),
      .za_waitrequest (sdram_0_s1_waitrequest),
      .zs_addr        (zs_addr_from_the_sdram_0),
      .zs_ba          (zs_ba_from_the_sdram_0),
      .zs_cas_n       (zs_cas_n_from_the_sdram_0),
      .zs_cke         (zs_cke_from_the_sdram_0),
      .zs_cs_n        (zs_cs_n_from_the_sdram_0),
      .zs_dq          (zs_dq_to_and_from_the_sdram_0),
      .zs_dqm         (zs_dqm_from_the_sdram_0),
      .zs_ras_n       (zs_ras_n_from_the_sdram_0),
      .zs_we_n        (zs_we_n_from_the_sdram_0)
    );

  sram_0_avalon_sram_slave_arbitrator the_sram_0_avalon_sram_slave
    (
      .clk                                                                                                      (sys_clk),
      .cpu_0_data_master_address_to_slave                                                                       (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                                                             (cpu_0_data_master_byteenable),
      .cpu_0_data_master_byteenable_sram_0_avalon_sram_slave                                                    (cpu_0_data_master_byteenable_sram_0_avalon_sram_slave),
      .cpu_0_data_master_dbs_address                                                                            (cpu_0_data_master_dbs_address),
      .cpu_0_data_master_dbs_write_16                                                                           (cpu_0_data_master_dbs_write_16),
      .cpu_0_data_master_granted_sram_0_avalon_sram_slave                                                       (cpu_0_data_master_granted_sram_0_avalon_sram_slave),
      .cpu_0_data_master_latency_counter                                                                        (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave                                             (cpu_0_data_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_0_data_master_read                                                                                   (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave                                               (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register                                (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_requests_sram_0_avalon_sram_slave                                                      (cpu_0_data_master_requests_sram_0_avalon_sram_slave),
      .cpu_0_data_master_write                                                                                  (cpu_0_data_master_write),
      .cpu_1_data_master_address_to_slave                                                                       (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_byteenable                                                                             (cpu_1_data_master_byteenable),
      .cpu_1_data_master_byteenable_sram_0_avalon_sram_slave                                                    (cpu_1_data_master_byteenable_sram_0_avalon_sram_slave),
      .cpu_1_data_master_dbs_address                                                                            (cpu_1_data_master_dbs_address),
      .cpu_1_data_master_dbs_write_16                                                                           (cpu_1_data_master_dbs_write_16),
      .cpu_1_data_master_granted_sram_0_avalon_sram_slave                                                       (cpu_1_data_master_granted_sram_0_avalon_sram_slave),
      .cpu_1_data_master_latency_counter                                                                        (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave                                             (cpu_1_data_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_1_data_master_read                                                                                   (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave                                               (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register                                (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_requests_sram_0_avalon_sram_slave                                                      (cpu_1_data_master_requests_sram_0_avalon_sram_slave),
      .cpu_1_data_master_write                                                                                  (cpu_1_data_master_write),
      .cpu_1_instruction_master_address_to_slave                                                                (cpu_1_instruction_master_address_to_slave),
      .cpu_1_instruction_master_dbs_address                                                                     (cpu_1_instruction_master_dbs_address),
      .cpu_1_instruction_master_granted_sram_0_avalon_sram_slave                                                (cpu_1_instruction_master_granted_sram_0_avalon_sram_slave),
      .cpu_1_instruction_master_latency_counter                                                                 (cpu_1_instruction_master_latency_counter),
      .cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave                                      (cpu_1_instruction_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_1_instruction_master_read                                                                            (cpu_1_instruction_master_read),
      .cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave                                        (cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register                         (cpu_1_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_instruction_master_requests_sram_0_avalon_sram_slave                                               (cpu_1_instruction_master_requests_sram_0_avalon_sram_slave),
      .cpu_2_data_master_address_to_slave                                                                       (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_byteenable                                                                             (cpu_2_data_master_byteenable),
      .cpu_2_data_master_byteenable_sram_0_avalon_sram_slave                                                    (cpu_2_data_master_byteenable_sram_0_avalon_sram_slave),
      .cpu_2_data_master_dbs_address                                                                            (cpu_2_data_master_dbs_address),
      .cpu_2_data_master_dbs_write_16                                                                           (cpu_2_data_master_dbs_write_16),
      .cpu_2_data_master_granted_sram_0_avalon_sram_slave                                                       (cpu_2_data_master_granted_sram_0_avalon_sram_slave),
      .cpu_2_data_master_latency_counter                                                                        (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave                                             (cpu_2_data_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_2_data_master_read                                                                                   (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave                                               (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register                                (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_requests_sram_0_avalon_sram_slave                                                      (cpu_2_data_master_requests_sram_0_avalon_sram_slave),
      .cpu_2_data_master_write                                                                                  (cpu_2_data_master_write),
      .cpu_2_instruction_master_address_to_slave                                                                (cpu_2_instruction_master_address_to_slave),
      .cpu_2_instruction_master_dbs_address                                                                     (cpu_2_instruction_master_dbs_address),
      .cpu_2_instruction_master_granted_sram_0_avalon_sram_slave                                                (cpu_2_instruction_master_granted_sram_0_avalon_sram_slave),
      .cpu_2_instruction_master_latency_counter                                                                 (cpu_2_instruction_master_latency_counter),
      .cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave                                      (cpu_2_instruction_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_2_instruction_master_read                                                                            (cpu_2_instruction_master_read),
      .cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave                                        (cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register                         (cpu_2_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_instruction_master_requests_sram_0_avalon_sram_slave                                               (cpu_2_instruction_master_requests_sram_0_avalon_sram_slave),
      .cpu_3_data_master_address_to_slave                                                                       (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_byteenable                                                                             (cpu_3_data_master_byteenable),
      .cpu_3_data_master_byteenable_sram_0_avalon_sram_slave                                                    (cpu_3_data_master_byteenable_sram_0_avalon_sram_slave),
      .cpu_3_data_master_dbs_address                                                                            (cpu_3_data_master_dbs_address),
      .cpu_3_data_master_dbs_write_16                                                                           (cpu_3_data_master_dbs_write_16),
      .cpu_3_data_master_granted_sram_0_avalon_sram_slave                                                       (cpu_3_data_master_granted_sram_0_avalon_sram_slave),
      .cpu_3_data_master_latency_counter                                                                        (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave                                             (cpu_3_data_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_3_data_master_read                                                                                   (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave                                               (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register                                (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_requests_sram_0_avalon_sram_slave                                                      (cpu_3_data_master_requests_sram_0_avalon_sram_slave),
      .cpu_3_data_master_write                                                                                  (cpu_3_data_master_write),
      .cpu_3_instruction_master_address_to_slave                                                                (cpu_3_instruction_master_address_to_slave),
      .cpu_3_instruction_master_dbs_address                                                                     (cpu_3_instruction_master_dbs_address),
      .cpu_3_instruction_master_granted_sram_0_avalon_sram_slave                                                (cpu_3_instruction_master_granted_sram_0_avalon_sram_slave),
      .cpu_3_instruction_master_latency_counter                                                                 (cpu_3_instruction_master_latency_counter),
      .cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave                                      (cpu_3_instruction_master_qualified_request_sram_0_avalon_sram_slave),
      .cpu_3_instruction_master_read                                                                            (cpu_3_instruction_master_read),
      .cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave                                        (cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave),
      .cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register                         (cpu_3_instruction_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_instruction_master_requests_sram_0_avalon_sram_slave                                               (cpu_3_instruction_master_requests_sram_0_avalon_sram_slave),
      .d1_sram_0_avalon_sram_slave_end_xfer                                                                     (d1_sram_0_avalon_sram_slave_end_xfer),
      .reset_n                                                                                                  (sys_clk_reset_n),
      .sram_0_avalon_sram_slave_address                                                                         (sram_0_avalon_sram_slave_address),
      .sram_0_avalon_sram_slave_byteenable                                                                      (sram_0_avalon_sram_slave_byteenable),
      .sram_0_avalon_sram_slave_read                                                                            (sram_0_avalon_sram_slave_read),
      .sram_0_avalon_sram_slave_readdata                                                                        (sram_0_avalon_sram_slave_readdata),
      .sram_0_avalon_sram_slave_readdata_from_sa                                                                (sram_0_avalon_sram_slave_readdata_from_sa),
      .sram_0_avalon_sram_slave_readdatavalid                                                                   (sram_0_avalon_sram_slave_readdatavalid),
      .sram_0_avalon_sram_slave_reset                                                                           (sram_0_avalon_sram_slave_reset),
      .sram_0_avalon_sram_slave_write                                                                           (sram_0_avalon_sram_slave_write),
      .sram_0_avalon_sram_slave_writedata                                                                       (sram_0_avalon_sram_slave_writedata),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave                                        (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock                                             (video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address                                             (video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave                        (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter                                         (video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave              (video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_read                                                    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave                (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave                       (video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave)
    );

  sram_0 the_sram_0
    (
      .SRAM_ADDR     (SRAM_ADDR_from_the_sram_0),
      .SRAM_CE_N     (SRAM_CE_N_from_the_sram_0),
      .SRAM_DQ       (SRAM_DQ_to_and_from_the_sram_0),
      .SRAM_LB_N     (SRAM_LB_N_from_the_sram_0),
      .SRAM_OE_N     (SRAM_OE_N_from_the_sram_0),
      .SRAM_UB_N     (SRAM_UB_N_from_the_sram_0),
      .SRAM_WE_N     (SRAM_WE_N_from_the_sram_0),
      .address       (sram_0_avalon_sram_slave_address),
      .byteenable    (sram_0_avalon_sram_slave_byteenable),
      .clk           (sys_clk),
      .read          (sram_0_avalon_sram_slave_read),
      .readdata      (sram_0_avalon_sram_slave_readdata),
      .readdatavalid (sram_0_avalon_sram_slave_readdatavalid),
      .reset         (sram_0_avalon_sram_slave_reset),
      .write         (sram_0_avalon_sram_slave_write),
      .writedata     (sram_0_avalon_sram_slave_writedata)
    );

  sysid_control_slave_arbitrator the_sysid_control_slave
    (
      .clk                                                                       (sys_clk),
      .cpu_0_data_master_address_to_slave                                        (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_sysid_control_slave                             (cpu_0_data_master_granted_sysid_control_slave),
      .cpu_0_data_master_latency_counter                                         (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_sysid_control_slave                   (cpu_0_data_master_qualified_request_sysid_control_slave),
      .cpu_0_data_master_read                                                    (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_read_data_valid_sysid_control_slave                     (cpu_0_data_master_read_data_valid_sysid_control_slave),
      .cpu_0_data_master_requests_sysid_control_slave                            (cpu_0_data_master_requests_sysid_control_slave),
      .cpu_0_data_master_write                                                   (cpu_0_data_master_write),
      .cpu_1_data_master_address_to_slave                                        (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_granted_sysid_control_slave                             (cpu_1_data_master_granted_sysid_control_slave),
      .cpu_1_data_master_latency_counter                                         (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_sysid_control_slave                   (cpu_1_data_master_qualified_request_sysid_control_slave),
      .cpu_1_data_master_read                                                    (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_read_data_valid_sysid_control_slave                     (cpu_1_data_master_read_data_valid_sysid_control_slave),
      .cpu_1_data_master_requests_sysid_control_slave                            (cpu_1_data_master_requests_sysid_control_slave),
      .cpu_1_data_master_write                                                   (cpu_1_data_master_write),
      .cpu_2_data_master_address_to_slave                                        (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_granted_sysid_control_slave                             (cpu_2_data_master_granted_sysid_control_slave),
      .cpu_2_data_master_latency_counter                                         (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_sysid_control_slave                   (cpu_2_data_master_qualified_request_sysid_control_slave),
      .cpu_2_data_master_read                                                    (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_read_data_valid_sysid_control_slave                     (cpu_2_data_master_read_data_valid_sysid_control_slave),
      .cpu_2_data_master_requests_sysid_control_slave                            (cpu_2_data_master_requests_sysid_control_slave),
      .cpu_2_data_master_write                                                   (cpu_2_data_master_write),
      .cpu_3_data_master_address_to_slave                                        (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_granted_sysid_control_slave                             (cpu_3_data_master_granted_sysid_control_slave),
      .cpu_3_data_master_latency_counter                                         (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_sysid_control_slave                   (cpu_3_data_master_qualified_request_sysid_control_slave),
      .cpu_3_data_master_read                                                    (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_read_data_valid_sysid_control_slave                     (cpu_3_data_master_read_data_valid_sysid_control_slave),
      .cpu_3_data_master_requests_sysid_control_slave                            (cpu_3_data_master_requests_sysid_control_slave),
      .cpu_3_data_master_write                                                   (cpu_3_data_master_write),
      .d1_sysid_control_slave_end_xfer                                           (d1_sysid_control_slave_end_xfer),
      .reset_n                                                                   (sys_clk_reset_n),
      .sysid_control_slave_address                                               (sysid_control_slave_address),
      .sysid_control_slave_readdata                                              (sysid_control_slave_readdata),
      .sysid_control_slave_readdata_from_sa                                      (sysid_control_slave_readdata_from_sa),
      .sysid_control_slave_reset_n                                               (sysid_control_slave_reset_n)
    );

  sysid the_sysid
    (
      .address  (sysid_control_slave_address),
      .clock    (sysid_control_slave_clock),
      .readdata (sysid_control_slave_readdata),
      .reset_n  (sysid_control_slave_reset_n)
    );

  video_dual_clock_buffer_0_avalon_dc_buffer_sink_arbitrator the_video_dual_clock_buffer_0_avalon_dc_buffer_sink
    (
      .clk                                                           (sys_clk),
      .reset_n                                                       (sys_clk_reset_n),
      .video_dual_clock_buffer_0_avalon_dc_buffer_sink_data          (video_dual_clock_buffer_0_avalon_dc_buffer_sink_data),
      .video_dual_clock_buffer_0_avalon_dc_buffer_sink_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_sink_endofpacket),
      .video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready),
      .video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa (video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa),
      .video_dual_clock_buffer_0_avalon_dc_buffer_sink_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_sink_startofpacket),
      .video_dual_clock_buffer_0_avalon_dc_buffer_sink_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_sink_valid),
      .video_scaler_0_avalon_scaler_source_data                      (video_scaler_0_avalon_scaler_source_data),
      .video_scaler_0_avalon_scaler_source_endofpacket               (video_scaler_0_avalon_scaler_source_endofpacket),
      .video_scaler_0_avalon_scaler_source_startofpacket             (video_scaler_0_avalon_scaler_source_startofpacket),
      .video_scaler_0_avalon_scaler_source_valid                     (video_scaler_0_avalon_scaler_source_valid)
    );

  video_dual_clock_buffer_0_avalon_dc_buffer_source_arbitrator the_video_dual_clock_buffer_0_avalon_dc_buffer_source
    (
      .clk                                                             (vga_clock),
      .reset_n                                                         (vga_clock_reset_n),
      .video_dual_clock_buffer_0_avalon_dc_buffer_source_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),
      .video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),
      .video_dual_clock_buffer_0_avalon_dc_buffer_source_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),
      .video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket),
      .video_dual_clock_buffer_0_avalon_dc_buffer_source_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),
      .video_vga_controller_0_avalon_vga_sink_ready_from_sa            (video_vga_controller_0_avalon_vga_sink_ready_from_sa)
    );

  video_dual_clock_buffer_0 the_video_dual_clock_buffer_0
    (
      .clk_stream_in            (sys_clk),
      .clk_stream_out           (vga_clock),
      .stream_in_data           (video_dual_clock_buffer_0_avalon_dc_buffer_sink_data),
      .stream_in_endofpacket    (video_dual_clock_buffer_0_avalon_dc_buffer_sink_endofpacket),
      .stream_in_ready          (video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready),
      .stream_in_startofpacket  (video_dual_clock_buffer_0_avalon_dc_buffer_sink_startofpacket),
      .stream_in_valid          (video_dual_clock_buffer_0_avalon_dc_buffer_sink_valid),
      .stream_out_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),
      .stream_out_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),
      .stream_out_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),
      .stream_out_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket),
      .stream_out_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid)
    );

  video_pixel_buffer_dma_0_avalon_control_slave_arbitrator the_video_pixel_buffer_dma_0_avalon_control_slave
    (
      .clk                                                                               (sys_clk),
      .cpu_0_data_master_address_to_slave                                                (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                                      (cpu_0_data_master_byteenable),
      .cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave           (cpu_0_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_0_data_master_latency_counter                                                 (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave (cpu_0_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_0_data_master_read                                                            (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register         (cpu_0_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave   (cpu_0_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave          (cpu_0_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_0_data_master_write                                                           (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                                       (cpu_0_data_master_writedata),
      .cpu_1_data_master_address_to_slave                                                (cpu_1_data_master_address_to_slave),
      .cpu_1_data_master_byteenable                                                      (cpu_1_data_master_byteenable),
      .cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave           (cpu_1_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_1_data_master_latency_counter                                                 (cpu_1_data_master_latency_counter),
      .cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave (cpu_1_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_1_data_master_read                                                            (cpu_1_data_master_read),
      .cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register         (cpu_1_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave   (cpu_1_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave          (cpu_1_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_1_data_master_write                                                           (cpu_1_data_master_write),
      .cpu_1_data_master_writedata                                                       (cpu_1_data_master_writedata),
      .cpu_2_data_master_address_to_slave                                                (cpu_2_data_master_address_to_slave),
      .cpu_2_data_master_byteenable                                                      (cpu_2_data_master_byteenable),
      .cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave           (cpu_2_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_2_data_master_latency_counter                                                 (cpu_2_data_master_latency_counter),
      .cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave (cpu_2_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_2_data_master_read                                                            (cpu_2_data_master_read),
      .cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register         (cpu_2_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave   (cpu_2_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave          (cpu_2_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_2_data_master_write                                                           (cpu_2_data_master_write),
      .cpu_2_data_master_writedata                                                       (cpu_2_data_master_writedata),
      .cpu_3_data_master_address_to_slave                                                (cpu_3_data_master_address_to_slave),
      .cpu_3_data_master_byteenable                                                      (cpu_3_data_master_byteenable),
      .cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave           (cpu_3_data_master_granted_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_3_data_master_latency_counter                                                 (cpu_3_data_master_latency_counter),
      .cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave (cpu_3_data_master_qualified_request_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_3_data_master_read                                                            (cpu_3_data_master_read),
      .cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register         (cpu_3_data_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave   (cpu_3_data_master_read_data_valid_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave          (cpu_3_data_master_requests_video_pixel_buffer_dma_0_avalon_control_slave),
      .cpu_3_data_master_write                                                           (cpu_3_data_master_write),
      .cpu_3_data_master_writedata                                                       (cpu_3_data_master_writedata),
      .d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer                         (d1_video_pixel_buffer_dma_0_avalon_control_slave_end_xfer),
      .reset_n                                                                           (sys_clk_reset_n),
      .video_pixel_buffer_dma_0_avalon_control_slave_address                             (video_pixel_buffer_dma_0_avalon_control_slave_address),
      .video_pixel_buffer_dma_0_avalon_control_slave_byteenable                          (video_pixel_buffer_dma_0_avalon_control_slave_byteenable),
      .video_pixel_buffer_dma_0_avalon_control_slave_read                                (video_pixel_buffer_dma_0_avalon_control_slave_read),
      .video_pixel_buffer_dma_0_avalon_control_slave_readdata                            (video_pixel_buffer_dma_0_avalon_control_slave_readdata),
      .video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa                    (video_pixel_buffer_dma_0_avalon_control_slave_readdata_from_sa),
      .video_pixel_buffer_dma_0_avalon_control_slave_write                               (video_pixel_buffer_dma_0_avalon_control_slave_write),
      .video_pixel_buffer_dma_0_avalon_control_slave_writedata                           (video_pixel_buffer_dma_0_avalon_control_slave_writedata)
    );

  video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbitrator the_video_pixel_buffer_dma_0_avalon_pixel_dma_master
    (
      .clk                                                                                                      (sys_clk),
      .d1_sram_0_avalon_sram_slave_end_xfer                                                                     (d1_sram_0_avalon_sram_slave_end_xfer),
      .reset_n                                                                                                  (sys_clk_reset_n),
      .sram_0_avalon_sram_slave_readdata_from_sa                                                                (sram_0_avalon_sram_slave_readdata_from_sa),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_address                                                 (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave                                        (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address_to_slave),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address                                             (video_pixel_buffer_dma_0_avalon_pixel_dma_master_dbs_address),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave                        (video_pixel_buffer_dma_0_avalon_pixel_dma_master_granted_sram_0_avalon_sram_slave),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter                                         (video_pixel_buffer_dma_0_avalon_pixel_dma_master_latency_counter),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave              (video_pixel_buffer_dma_0_avalon_pixel_dma_master_qualified_request_sram_0_avalon_sram_slave),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_read                                                    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave                (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave_shift_register (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read_data_valid_sram_0_avalon_sram_slave_shift_register),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata                                                (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid                                           (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave                       (video_pixel_buffer_dma_0_avalon_pixel_dma_master_requests_sram_0_avalon_sram_slave),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_reset                                                   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_reset),
      .video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest                                             (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest)
    );

  video_pixel_buffer_dma_0_avalon_pixel_source_arbitrator the_video_pixel_buffer_dma_0_avalon_pixel_source
    (
      .clk                                                        (sys_clk),
      .reset_n                                                    (sys_clk_reset_n),
      .video_pixel_buffer_dma_0_avalon_pixel_source_data          (video_pixel_buffer_dma_0_avalon_pixel_source_data),
      .video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket   (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),
      .video_pixel_buffer_dma_0_avalon_pixel_source_ready         (video_pixel_buffer_dma_0_avalon_pixel_source_ready),
      .video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket),
      .video_pixel_buffer_dma_0_avalon_pixel_source_valid         (video_pixel_buffer_dma_0_avalon_pixel_source_valid),
      .video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa        (video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa)
    );

  video_pixel_buffer_dma_0 the_video_pixel_buffer_dma_0
    (
      .clk                  (sys_clk),
      .master_address       (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),
      .master_arbiterlock   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_arbiterlock),
      .master_read          (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),
      .master_readdata      (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),
      .master_readdatavalid (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),
      .master_waitrequest   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),
      .reset                (video_pixel_buffer_dma_0_avalon_pixel_dma_master_reset),
      .slave_address        (video_pixel_buffer_dma_0_avalon_control_slave_address),
      .slave_byteenable     (video_pixel_buffer_dma_0_avalon_control_slave_byteenable),
      .slave_read           (video_pixel_buffer_dma_0_avalon_control_slave_read),
      .slave_readdata       (video_pixel_buffer_dma_0_avalon_control_slave_readdata),
      .slave_write          (video_pixel_buffer_dma_0_avalon_control_slave_write),
      .slave_writedata      (video_pixel_buffer_dma_0_avalon_control_slave_writedata),
      .stream_data          (video_pixel_buffer_dma_0_avalon_pixel_source_data),
      .stream_endofpacket   (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),
      .stream_ready         (video_pixel_buffer_dma_0_avalon_pixel_source_ready),
      .stream_startofpacket (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket),
      .stream_valid         (video_pixel_buffer_dma_0_avalon_pixel_source_valid)
    );

  video_rgb_resampler_0_avalon_rgb_sink_arbitrator the_video_rgb_resampler_0_avalon_rgb_sink
    (
      .clk                                                        (sys_clk),
      .reset_n                                                    (sys_clk_reset_n),
      .video_pixel_buffer_dma_0_avalon_pixel_source_data          (video_pixel_buffer_dma_0_avalon_pixel_source_data),
      .video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket   (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),
      .video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket),
      .video_pixel_buffer_dma_0_avalon_pixel_source_valid         (video_pixel_buffer_dma_0_avalon_pixel_source_valid),
      .video_rgb_resampler_0_avalon_rgb_sink_data                 (video_rgb_resampler_0_avalon_rgb_sink_data),
      .video_rgb_resampler_0_avalon_rgb_sink_endofpacket          (video_rgb_resampler_0_avalon_rgb_sink_endofpacket),
      .video_rgb_resampler_0_avalon_rgb_sink_ready                (video_rgb_resampler_0_avalon_rgb_sink_ready),
      .video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa        (video_rgb_resampler_0_avalon_rgb_sink_ready_from_sa),
      .video_rgb_resampler_0_avalon_rgb_sink_reset                (video_rgb_resampler_0_avalon_rgb_sink_reset),
      .video_rgb_resampler_0_avalon_rgb_sink_startofpacket        (video_rgb_resampler_0_avalon_rgb_sink_startofpacket),
      .video_rgb_resampler_0_avalon_rgb_sink_valid                (video_rgb_resampler_0_avalon_rgb_sink_valid)
    );

  video_rgb_resampler_0_avalon_rgb_source_arbitrator the_video_rgb_resampler_0_avalon_rgb_source
    (
      .clk                                                   (sys_clk),
      .reset_n                                               (sys_clk_reset_n),
      .video_rgb_resampler_0_avalon_rgb_source_data          (video_rgb_resampler_0_avalon_rgb_source_data),
      .video_rgb_resampler_0_avalon_rgb_source_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),
      .video_rgb_resampler_0_avalon_rgb_source_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),
      .video_rgb_resampler_0_avalon_rgb_source_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),
      .video_rgb_resampler_0_avalon_rgb_source_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),
      .video_scaler_0_avalon_scaler_sink_ready_from_sa       (video_scaler_0_avalon_scaler_sink_ready_from_sa)
    );

  video_rgb_resampler_0 the_video_rgb_resampler_0
    (
      .clk                      (sys_clk),
      .reset                    (video_rgb_resampler_0_avalon_rgb_sink_reset),
      .stream_in_data           (video_rgb_resampler_0_avalon_rgb_sink_data),
      .stream_in_endofpacket    (video_rgb_resampler_0_avalon_rgb_sink_endofpacket),
      .stream_in_ready          (video_rgb_resampler_0_avalon_rgb_sink_ready),
      .stream_in_startofpacket  (video_rgb_resampler_0_avalon_rgb_sink_startofpacket),
      .stream_in_valid          (video_rgb_resampler_0_avalon_rgb_sink_valid),
      .stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data),
      .stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),
      .stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),
      .stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),
      .stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid)
    );

  video_scaler_0_avalon_scaler_sink_arbitrator the_video_scaler_0_avalon_scaler_sink
    (
      .clk                                                   (sys_clk),
      .reset_n                                               (sys_clk_reset_n),
      .video_rgb_resampler_0_avalon_rgb_source_data          (video_rgb_resampler_0_avalon_rgb_source_data),
      .video_rgb_resampler_0_avalon_rgb_source_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),
      .video_rgb_resampler_0_avalon_rgb_source_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),
      .video_rgb_resampler_0_avalon_rgb_source_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),
      .video_scaler_0_avalon_scaler_sink_data                (video_scaler_0_avalon_scaler_sink_data),
      .video_scaler_0_avalon_scaler_sink_endofpacket         (video_scaler_0_avalon_scaler_sink_endofpacket),
      .video_scaler_0_avalon_scaler_sink_ready               (video_scaler_0_avalon_scaler_sink_ready),
      .video_scaler_0_avalon_scaler_sink_ready_from_sa       (video_scaler_0_avalon_scaler_sink_ready_from_sa),
      .video_scaler_0_avalon_scaler_sink_reset               (video_scaler_0_avalon_scaler_sink_reset),
      .video_scaler_0_avalon_scaler_sink_startofpacket       (video_scaler_0_avalon_scaler_sink_startofpacket),
      .video_scaler_0_avalon_scaler_sink_valid               (video_scaler_0_avalon_scaler_sink_valid)
    );

  video_scaler_0_avalon_scaler_source_arbitrator the_video_scaler_0_avalon_scaler_source
    (
      .clk                                                           (sys_clk),
      .reset_n                                                       (sys_clk_reset_n),
      .video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa (video_dual_clock_buffer_0_avalon_dc_buffer_sink_ready_from_sa),
      .video_scaler_0_avalon_scaler_source_data                      (video_scaler_0_avalon_scaler_source_data),
      .video_scaler_0_avalon_scaler_source_endofpacket               (video_scaler_0_avalon_scaler_source_endofpacket),
      .video_scaler_0_avalon_scaler_source_ready                     (video_scaler_0_avalon_scaler_source_ready),
      .video_scaler_0_avalon_scaler_source_startofpacket             (video_scaler_0_avalon_scaler_source_startofpacket),
      .video_scaler_0_avalon_scaler_source_valid                     (video_scaler_0_avalon_scaler_source_valid)
    );

  video_scaler_0 the_video_scaler_0
    (
      .clk                      (sys_clk),
      .reset                    (video_scaler_0_avalon_scaler_sink_reset),
      .stream_in_data           (video_scaler_0_avalon_scaler_sink_data),
      .stream_in_endofpacket    (video_scaler_0_avalon_scaler_sink_endofpacket),
      .stream_in_ready          (video_scaler_0_avalon_scaler_sink_ready),
      .stream_in_startofpacket  (video_scaler_0_avalon_scaler_sink_startofpacket),
      .stream_in_valid          (video_scaler_0_avalon_scaler_sink_valid),
      .stream_out_data          (video_scaler_0_avalon_scaler_source_data),
      .stream_out_endofpacket   (video_scaler_0_avalon_scaler_source_endofpacket),
      .stream_out_ready         (video_scaler_0_avalon_scaler_source_ready),
      .stream_out_startofpacket (video_scaler_0_avalon_scaler_source_startofpacket),
      .stream_out_valid         (video_scaler_0_avalon_scaler_source_valid)
    );

  video_vga_controller_0_avalon_vga_sink_arbitrator the_video_vga_controller_0_avalon_vga_sink
    (
      .clk                                                             (vga_clock),
      .reset_n                                                         (vga_clock_reset_n),
      .video_dual_clock_buffer_0_avalon_dc_buffer_source_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),
      .video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),
      .video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket),
      .video_dual_clock_buffer_0_avalon_dc_buffer_source_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),
      .video_vga_controller_0_avalon_vga_sink_data                     (video_vga_controller_0_avalon_vga_sink_data),
      .video_vga_controller_0_avalon_vga_sink_endofpacket              (video_vga_controller_0_avalon_vga_sink_endofpacket),
      .video_vga_controller_0_avalon_vga_sink_ready                    (video_vga_controller_0_avalon_vga_sink_ready),
      .video_vga_controller_0_avalon_vga_sink_ready_from_sa            (video_vga_controller_0_avalon_vga_sink_ready_from_sa),
      .video_vga_controller_0_avalon_vga_sink_reset                    (video_vga_controller_0_avalon_vga_sink_reset),
      .video_vga_controller_0_avalon_vga_sink_startofpacket            (video_vga_controller_0_avalon_vga_sink_startofpacket),
      .video_vga_controller_0_avalon_vga_sink_valid                    (video_vga_controller_0_avalon_vga_sink_valid)
    );

  video_vga_controller_0 the_video_vga_controller_0
    (
      .VGA_B         (VGA_B_from_the_video_vga_controller_0),
      .VGA_BLANK     (VGA_BLANK_from_the_video_vga_controller_0),
      .VGA_CLK       (VGA_CLK_from_the_video_vga_controller_0),
      .VGA_G         (VGA_G_from_the_video_vga_controller_0),
      .VGA_HS        (VGA_HS_from_the_video_vga_controller_0),
      .VGA_R         (VGA_R_from_the_video_vga_controller_0),
      .VGA_SYNC      (VGA_SYNC_from_the_video_vga_controller_0),
      .VGA_VS        (VGA_VS_from_the_video_vga_controller_0),
      .clk           (vga_clock),
      .data          (video_vga_controller_0_avalon_vga_sink_data),
      .endofpacket   (video_vga_controller_0_avalon_vga_sink_endofpacket),
      .ready         (video_vga_controller_0_avalon_vga_sink_ready),
      .reset         (video_vga_controller_0_avalon_vga_sink_reset),
      .startofpacket (video_vga_controller_0_avalon_vga_sink_startofpacket),
      .valid         (video_vga_controller_0_avalon_vga_sink_valid)
    );

  //reset is asserted asynchronously and deasserted synchronously
  nios_system_reset_clk_0_domain_synch_module nios_system_reset_clk_0_domain_synch
    (
      .clk      (clk_0),
      .data_in  (1'b1),
      .data_out (clk_0_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset sources mux, which is an e_mux
  assign reset_n_sources = ~(~reset_n |
    0 |
    0 |
    cpu_0_jtag_debug_module_resetrequest_from_sa |
    cpu_0_jtag_debug_module_resetrequest_from_sa |
    cpu_1_jtag_debug_module_resetrequest_from_sa |
    cpu_1_jtag_debug_module_resetrequest_from_sa |
    cpu_2_jtag_debug_module_resetrequest_from_sa |
    cpu_2_jtag_debug_module_resetrequest_from_sa |
    cpu_3_jtag_debug_module_resetrequest_from_sa |
    cpu_3_jtag_debug_module_resetrequest_from_sa |
    0 |
    0);

  //reset is asserted asynchronously and deasserted synchronously
  nios_system_reset_sys_clk_domain_synch_module nios_system_reset_sys_clk_domain_synch
    (
      .clk      (sys_clk),
      .data_in  (1'b1),
      .data_out (sys_clk_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset is asserted asynchronously and deasserted synchronously
  nios_system_reset_sdram_clk_domain_synch_module nios_system_reset_sdram_clk_domain_synch
    (
      .clk      (sdram_clk),
      .data_in  (1'b1),
      .data_out (sdram_clk_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset is asserted asynchronously and deasserted synchronously
  nios_system_reset_vga_clock_domain_synch_module nios_system_reset_vga_clock_domain_synch
    (
      .clk      (vga_clock),
      .data_in  (1'b1),
      .data_out (vga_clock_reset_n),
      .reset_n  (reset_n_sources)
    );

  //nios_system_clock_0_in_writedata of type writedata does not connect to anything so wire it to default (0)
  assign nios_system_clock_0_in_writedata = 0;

  //nios_system_clock_0_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_0_out_endofpacket = 0;

  //nios_system_clock_10_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_10_out_endofpacket = 0;

  //nios_system_clock_11_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_11_out_endofpacket = 0;

  //nios_system_clock_1_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_1_out_endofpacket = 0;

  //nios_system_clock_2_in_writedata of type writedata does not connect to anything so wire it to default (0)
  assign nios_system_clock_2_in_writedata = 0;

  //nios_system_clock_2_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_2_out_endofpacket = 0;

  //nios_system_clock_3_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_3_out_endofpacket = 0;

  //nios_system_clock_4_in_writedata of type writedata does not connect to anything so wire it to default (0)
  assign nios_system_clock_4_in_writedata = 0;

  //nios_system_clock_4_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_4_out_endofpacket = 0;

  //nios_system_clock_5_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_5_out_endofpacket = 0;

  //nios_system_clock_6_in_writedata of type writedata does not connect to anything so wire it to default (0)
  assign nios_system_clock_6_in_writedata = 0;

  //nios_system_clock_6_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_6_out_endofpacket = 0;

  //nios_system_clock_7_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_7_out_endofpacket = 0;

  //nios_system_clock_8_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_8_out_endofpacket = 0;

  //nios_system_clock_9_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign nios_system_clock_9_out_endofpacket = 0;

  //sysid_control_slave_clock of type clock does not connect to anything so wire it to default (0)
  assign sysid_control_slave_clock = 0;


endmodule


//synthesis translate_off



// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE

// AND HERE WILL BE PRESERVED </ALTERA_NOTE>


// If user logic components use Altsync_Ram with convert_hex2ver.dll,
// set USE_convert_hex2ver in the user comments section above

// `ifdef USE_convert_hex2ver
// `else
// `define NO_PLI 1
// `endif

`include "/usr/local/3rdparty/altera/quartus12/quartus/eda/sim_lib/altera_mf.v"
`include "/usr/local/3rdparty/altera/quartus12/quartus/eda/sim_lib/220model.v"
`include "/usr/local/3rdparty/altera/quartus12/quartus/eda/sim_lib/sgate.v"
`include "sram_0.v"
`include "/usr/local/3rdparty/altera/quartus12/ip/altera/nios2_ip/altera_nios_custom_instr_floating_point_qsys/fpoint_wrapper.v"
`include "/usr/local/3rdparty/altera/quartus12/ip/altera/nios2_ip/altera_nios_custom_instr_floating_point_qsys/fpoint_qsys.v"
`include "/usr/local/3rdparty/altera/quartus12/ip/altera/nios2_ip/altera_nios_custom_instr_floating_point_qsys/fpoint_hw_qsys.v"
`include "cpu_2_altera_nios_custom_instr_floating_point_inst.v"
`include "clocks_0.v"
`include "video_dual_clock_buffer_0.v"
`include "video_rgb_resampler_0.v"
`include "video_scaler_0.v"
`include "video_vga_controller_0.v"
`include "cpu_3_altera_nios_custom_instr_floating_point_inst.v"
`include "cpu_1_altera_nios_custom_instr_floating_point_inst.v"
`include "cpu_0_altera_nios_custom_instr_floating_point_inst.v"
`include "video_pixel_buffer_dma_0.v"
`include "jtag_uart_1.v"
`include "nios_system_clock_8.v"
`include "cpu_2_test_bench.v"
`include "cpu_2_mult_cell.v"
`include "cpu_2_oci_test_bench.v"
`include "cpu_2_jtag_debug_module_tck.v"
`include "cpu_2_jtag_debug_module_sysclk.v"
`include "cpu_2_jtag_debug_module_wrapper.v"
`include "cpu_2.v"
`include "onchip_memory2_1.v"
`include "nios_system_clock_1.v"
`include "sysid.v"
`include "cpu_0_test_bench.v"
`include "cpu_0_mult_cell.v"
`include "cpu_0_oci_test_bench.v"
`include "cpu_0_jtag_debug_module_tck.v"
`include "cpu_0_jtag_debug_module_sysclk.v"
`include "cpu_0_jtag_debug_module_wrapper.v"
`include "cpu_0.v"
`include "nios_system_clock_5.v"
`include "nios_system_clock_4.v"
`include "jtag_uart_0.v"
`include "onchip_memory2_0.v"
`include "cpu_1_test_bench.v"
`include "cpu_1_mult_cell.v"
`include "cpu_1_oci_test_bench.v"
`include "cpu_1_jtag_debug_module_tck.v"
`include "cpu_1_jtag_debug_module_sysclk.v"
`include "cpu_1_jtag_debug_module_wrapper.v"
`include "cpu_1.v"
`include "sdram_0.v"
`include "nios_system_clock_9.v"
`include "nios_system_clock_2.v"
`include "cpu_3_test_bench.v"
`include "cpu_3_mult_cell.v"
`include "cpu_3_oci_test_bench.v"
`include "cpu_3_jtag_debug_module_tck.v"
`include "cpu_3_jtag_debug_module_sysclk.v"
`include "cpu_3_jtag_debug_module_wrapper.v"
`include "cpu_3.v"
`include "jtag_uart_2.v"
`include "onchip_memory2_3.v"
`include "jtag_uart_3.v"
`include "nios_system_clock_0.v"
`include "mailbox_3.v"
`include "nios_system_clock_10.v"
`include "onchip_memory2_2.v"
`include "nios_system_clock_3.v"
`include "keys.v"
`include "mailbox_2.v"
`include "nios_system_clock_11.v"
`include "nios_system_clock_7.v"
`include "nios_system_clock_6.v"
`include "mailbox_1.v"
`include "performance_counter_0.v"
`include "mailbox_0.v"

`timescale 1ns / 1ps

module test_bench 
;


  wire    [ 17: 0] SRAM_ADDR_from_the_sram_0;
  wire             SRAM_CE_N_from_the_sram_0;
  wire    [ 15: 0] SRAM_DQ_to_and_from_the_sram_0;
  wire             SRAM_LB_N_from_the_sram_0;
  wire             SRAM_OE_N_from_the_sram_0;
  wire             SRAM_UB_N_from_the_sram_0;
  wire             SRAM_WE_N_from_the_sram_0;
  wire             VGA_BLANK_from_the_video_vga_controller_0;
  wire    [  9: 0] VGA_B_from_the_video_vga_controller_0;
  wire             VGA_CLK_from_the_video_vga_controller_0;
  wire    [  9: 0] VGA_G_from_the_video_vga_controller_0;
  wire             VGA_HS_from_the_video_vga_controller_0;
  wire    [  9: 0] VGA_R_from_the_video_vga_controller_0;
  wire             VGA_SYNC_from_the_video_vga_controller_0;
  wire             VGA_VS_from_the_video_vga_controller_0;
  wire             clk;
  reg              clk_0;
  wire    [  4: 0] cpu_0_custom_instruction_master_multi_a;
  wire    [  4: 0] cpu_0_custom_instruction_master_multi_b;
  wire    [  4: 0] cpu_0_custom_instruction_master_multi_c;
  wire             cpu_0_custom_instruction_master_multi_clk;
  wire             cpu_0_custom_instruction_master_multi_estatus;
  wire    [ 31: 0] cpu_0_custom_instruction_master_multi_ipending;
  wire             cpu_0_custom_instruction_master_multi_readra;
  wire             cpu_0_custom_instruction_master_multi_readrb;
  wire             cpu_0_custom_instruction_master_multi_reset;
  wire             cpu_0_custom_instruction_master_multi_status;
  wire             cpu_0_custom_instruction_master_multi_writerc;
  wire    [  4: 0] cpu_1_custom_instruction_master_multi_a;
  wire    [  4: 0] cpu_1_custom_instruction_master_multi_b;
  wire    [  4: 0] cpu_1_custom_instruction_master_multi_c;
  wire             cpu_1_custom_instruction_master_multi_clk;
  wire             cpu_1_custom_instruction_master_multi_estatus;
  wire    [ 31: 0] cpu_1_custom_instruction_master_multi_ipending;
  wire             cpu_1_custom_instruction_master_multi_readra;
  wire             cpu_1_custom_instruction_master_multi_readrb;
  wire             cpu_1_custom_instruction_master_multi_reset;
  wire             cpu_1_custom_instruction_master_multi_status;
  wire             cpu_1_custom_instruction_master_multi_writerc;
  wire    [  4: 0] cpu_2_custom_instruction_master_multi_a;
  wire    [  4: 0] cpu_2_custom_instruction_master_multi_b;
  wire    [  4: 0] cpu_2_custom_instruction_master_multi_c;
  wire             cpu_2_custom_instruction_master_multi_clk;
  wire             cpu_2_custom_instruction_master_multi_estatus;
  wire    [ 31: 0] cpu_2_custom_instruction_master_multi_ipending;
  wire             cpu_2_custom_instruction_master_multi_readra;
  wire             cpu_2_custom_instruction_master_multi_readrb;
  wire             cpu_2_custom_instruction_master_multi_reset;
  wire             cpu_2_custom_instruction_master_multi_status;
  wire             cpu_2_custom_instruction_master_multi_writerc;
  wire    [  4: 0] cpu_3_custom_instruction_master_multi_a;
  wire    [  4: 0] cpu_3_custom_instruction_master_multi_b;
  wire    [  4: 0] cpu_3_custom_instruction_master_multi_c;
  wire             cpu_3_custom_instruction_master_multi_clk;
  wire             cpu_3_custom_instruction_master_multi_estatus;
  wire    [ 31: 0] cpu_3_custom_instruction_master_multi_ipending;
  wire             cpu_3_custom_instruction_master_multi_readra;
  wire             cpu_3_custom_instruction_master_multi_readrb;
  wire             cpu_3_custom_instruction_master_multi_reset;
  wire             cpu_3_custom_instruction_master_multi_status;
  wire             cpu_3_custom_instruction_master_multi_writerc;
  wire    [  2: 0] in_port_to_the_keys;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_1_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_1_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_2_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_2_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_3_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_3_avalon_jtag_slave_readyfordata_from_sa;
  wire             nios_system_clock_0_in_endofpacket_from_sa;
  wire    [ 15: 0] nios_system_clock_0_in_writedata;
  wire             nios_system_clock_0_out_endofpacket;
  wire    [ 21: 0] nios_system_clock_0_out_nativeaddress;
  wire             nios_system_clock_10_in_endofpacket_from_sa;
  wire             nios_system_clock_10_out_endofpacket;
  wire             nios_system_clock_10_out_nativeaddress;
  wire             nios_system_clock_11_in_endofpacket_from_sa;
  wire             nios_system_clock_11_out_endofpacket;
  wire             nios_system_clock_11_out_nativeaddress;
  wire             nios_system_clock_1_in_endofpacket_from_sa;
  wire             nios_system_clock_1_out_endofpacket;
  wire    [ 21: 0] nios_system_clock_1_out_nativeaddress;
  wire             nios_system_clock_2_in_endofpacket_from_sa;
  wire    [ 15: 0] nios_system_clock_2_in_writedata;
  wire             nios_system_clock_2_out_endofpacket;
  wire    [ 21: 0] nios_system_clock_2_out_nativeaddress;
  wire             nios_system_clock_3_in_endofpacket_from_sa;
  wire             nios_system_clock_3_out_endofpacket;
  wire    [ 21: 0] nios_system_clock_3_out_nativeaddress;
  wire             nios_system_clock_4_in_endofpacket_from_sa;
  wire    [ 15: 0] nios_system_clock_4_in_writedata;
  wire             nios_system_clock_4_out_endofpacket;
  wire    [ 21: 0] nios_system_clock_4_out_nativeaddress;
  wire             nios_system_clock_5_in_endofpacket_from_sa;
  wire             nios_system_clock_5_out_endofpacket;
  wire    [ 21: 0] nios_system_clock_5_out_nativeaddress;
  wire             nios_system_clock_6_in_endofpacket_from_sa;
  wire    [ 15: 0] nios_system_clock_6_in_writedata;
  wire             nios_system_clock_6_out_endofpacket;
  wire    [ 21: 0] nios_system_clock_6_out_nativeaddress;
  wire             nios_system_clock_7_in_endofpacket_from_sa;
  wire             nios_system_clock_7_out_endofpacket;
  wire    [ 21: 0] nios_system_clock_7_out_nativeaddress;
  wire             nios_system_clock_8_in_endofpacket_from_sa;
  wire             nios_system_clock_8_out_endofpacket;
  wire             nios_system_clock_8_out_nativeaddress;
  wire             nios_system_clock_9_in_endofpacket_from_sa;
  wire             nios_system_clock_9_out_endofpacket;
  wire             nios_system_clock_9_out_nativeaddress;
  reg              reset_n;
  wire             sdram_clk;
  wire             sys_clk;
  wire             sysid_control_slave_clock;
  wire             vga_clock;
  wire    [ 11: 0] zs_addr_from_the_sdram_0;
  wire    [  1: 0] zs_ba_from_the_sdram_0;
  wire             zs_cas_n_from_the_sdram_0;
  wire             zs_cke_from_the_sdram_0;
  wire             zs_cs_n_from_the_sdram_0;
  wire    [ 15: 0] zs_dq_to_and_from_the_sdram_0;
  wire    [  1: 0] zs_dqm_from_the_sdram_0;
  wire             zs_ras_n_from_the_sdram_0;
  wire             zs_we_n_from_the_sdram_0;


// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
//  add your signals and additional architecture here
// AND HERE WILL BE PRESERVED </ALTERA_NOTE>

  //Set us up the Dut
  nios_system DUT
    (
      .SRAM_ADDR_from_the_sram_0                 (SRAM_ADDR_from_the_sram_0),
      .SRAM_CE_N_from_the_sram_0                 (SRAM_CE_N_from_the_sram_0),
      .SRAM_DQ_to_and_from_the_sram_0            (SRAM_DQ_to_and_from_the_sram_0),
      .SRAM_LB_N_from_the_sram_0                 (SRAM_LB_N_from_the_sram_0),
      .SRAM_OE_N_from_the_sram_0                 (SRAM_OE_N_from_the_sram_0),
      .SRAM_UB_N_from_the_sram_0                 (SRAM_UB_N_from_the_sram_0),
      .SRAM_WE_N_from_the_sram_0                 (SRAM_WE_N_from_the_sram_0),
      .VGA_BLANK_from_the_video_vga_controller_0 (VGA_BLANK_from_the_video_vga_controller_0),
      .VGA_B_from_the_video_vga_controller_0     (VGA_B_from_the_video_vga_controller_0),
      .VGA_CLK_from_the_video_vga_controller_0   (VGA_CLK_from_the_video_vga_controller_0),
      .VGA_G_from_the_video_vga_controller_0     (VGA_G_from_the_video_vga_controller_0),
      .VGA_HS_from_the_video_vga_controller_0    (VGA_HS_from_the_video_vga_controller_0),
      .VGA_R_from_the_video_vga_controller_0     (VGA_R_from_the_video_vga_controller_0),
      .VGA_SYNC_from_the_video_vga_controller_0  (VGA_SYNC_from_the_video_vga_controller_0),
      .VGA_VS_from_the_video_vga_controller_0    (VGA_VS_from_the_video_vga_controller_0),
      .clk_0                                     (clk_0),
      .in_port_to_the_keys                       (in_port_to_the_keys),
      .reset_n                                   (reset_n),
      .sdram_clk                                 (sdram_clk),
      .sys_clk                                   (sys_clk),
      .vga_clock                                 (vga_clock),
      .zs_addr_from_the_sdram_0                  (zs_addr_from_the_sdram_0),
      .zs_ba_from_the_sdram_0                    (zs_ba_from_the_sdram_0),
      .zs_cas_n_from_the_sdram_0                 (zs_cas_n_from_the_sdram_0),
      .zs_cke_from_the_sdram_0                   (zs_cke_from_the_sdram_0),
      .zs_cs_n_from_the_sdram_0                  (zs_cs_n_from_the_sdram_0),
      .zs_dq_to_and_from_the_sdram_0             (zs_dq_to_and_from_the_sdram_0),
      .zs_dqm_from_the_sdram_0                   (zs_dqm_from_the_sdram_0),
      .zs_ras_n_from_the_sdram_0                 (zs_ras_n_from_the_sdram_0),
      .zs_we_n_from_the_sdram_0                  (zs_we_n_from_the_sdram_0)
    );

  initial
    clk_0 = 1'b0;
  always
    #10 clk_0 <= ~clk_0;
  
  initial 
    begin
      reset_n <= 0;
      #200 reset_n <= 1;
    end

endmodule


//synthesis translate_on